module hanncoeffs4000(
	input wire [11:0]index,
	output reg signed [9:0]coeff
	);
	always @(index)
		case(index)
		12'd0: coeff = 10'sd0;
		12'd1: coeff = 10'sd0;
		12'd2: coeff = 10'sd0;
		12'd3: coeff = 10'sd0;
		12'd4: coeff = 10'sd0;
		12'd5: coeff = 10'sd0;
		12'd6: coeff = 10'sd0;
		12'd7: coeff = 10'sd0;
		12'd8: coeff = 10'sd0;
		12'd9: coeff = 10'sd0;
		12'd10: coeff = 10'sd0;
		12'd11: coeff = 10'sd0;
		12'd12: coeff = 10'sd0;
		12'd13: coeff = 10'sd0;
		12'd14: coeff = 10'sd0;
		12'd15: coeff = 10'sd0;
		12'd16: coeff = 10'sd0;
		12'd17: coeff = 10'sd0;
		12'd18: coeff = 10'sd0;
		12'd19: coeff = 10'sd0;
		12'd20: coeff = 10'sd0;
		12'd21: coeff = 10'sd0;
		12'd22: coeff = 10'sd0;
		12'd23: coeff = 10'sd0;
		12'd24: coeff = 10'sd0;
		12'd25: coeff = 10'sd0;
		12'd26: coeff = 10'sd0;
		12'd27: coeff = 10'sd0;
		12'd28: coeff = 10'sd0;
		12'd29: coeff = 10'sd1;
		12'd30: coeff = 10'sd1;
		12'd31: coeff = 10'sd1;
		12'd32: coeff = 10'sd1;
		12'd33: coeff = 10'sd1;
		12'd34: coeff = 10'sd1;
		12'd35: coeff = 10'sd1;
		12'd36: coeff = 10'sd1;
		12'd37: coeff = 10'sd1;
		12'd38: coeff = 10'sd1;
		12'd39: coeff = 10'sd1;
		12'd40: coeff = 10'sd1;
		12'd41: coeff = 10'sd1;
		12'd42: coeff = 10'sd1;
		12'd43: coeff = 10'sd1;
		12'd44: coeff = 10'sd1;
		12'd45: coeff = 10'sd1;
		12'd46: coeff = 10'sd1;
		12'd47: coeff = 10'sd1;
		12'd48: coeff = 10'sd1;
		12'd49: coeff = 10'sd2;
		12'd50: coeff = 10'sd2;
		12'd51: coeff = 10'sd2;
		12'd52: coeff = 10'sd2;
		12'd53: coeff = 10'sd2;
		12'd54: coeff = 10'sd2;
		12'd55: coeff = 10'sd2;
		12'd56: coeff = 10'sd2;
		12'd57: coeff = 10'sd2;
		12'd58: coeff = 10'sd2;
		12'd59: coeff = 10'sd2;
		12'd60: coeff = 10'sd2;
		12'd61: coeff = 10'sd2;
		12'd62: coeff = 10'sd2;
		12'd63: coeff = 10'sd3;
		12'd64: coeff = 10'sd3;
		12'd65: coeff = 10'sd3;
		12'd66: coeff = 10'sd3;
		12'd67: coeff = 10'sd3;
		12'd68: coeff = 10'sd3;
		12'd69: coeff = 10'sd3;
		12'd70: coeff = 10'sd3;
		12'd71: coeff = 10'sd3;
		12'd72: coeff = 10'sd3;
		12'd73: coeff = 10'sd3;
		12'd74: coeff = 10'sd3;
		12'd75: coeff = 10'sd4;
		12'd76: coeff = 10'sd4;
		12'd77: coeff = 10'sd4;
		12'd78: coeff = 10'sd4;
		12'd79: coeff = 10'sd4;
		12'd80: coeff = 10'sd4;
		12'd81: coeff = 10'sd4;
		12'd82: coeff = 10'sd4;
		12'd83: coeff = 10'sd4;
		12'd84: coeff = 10'sd4;
		12'd85: coeff = 10'sd5;
		12'd86: coeff = 10'sd5;
		12'd87: coeff = 10'sd5;
		12'd88: coeff = 10'sd5;
		12'd89: coeff = 10'sd5;
		12'd90: coeff = 10'sd5;
		12'd91: coeff = 10'sd5;
		12'd92: coeff = 10'sd5;
		12'd93: coeff = 10'sd5;
		12'd94: coeff = 10'sd6;
		12'd95: coeff = 10'sd6;
		12'd96: coeff = 10'sd6;
		12'd97: coeff = 10'sd6;
		12'd98: coeff = 10'sd6;
		12'd99: coeff = 10'sd6;
		12'd100: coeff = 10'sd6;
		12'd101: coeff = 10'sd6;
		12'd102: coeff = 10'sd7;
		12'd103: coeff = 10'sd7;
		12'd104: coeff = 10'sd7;
		12'd105: coeff = 10'sd7;
		12'd106: coeff = 10'sd7;
		12'd107: coeff = 10'sd7;
		12'd108: coeff = 10'sd7;
		12'd109: coeff = 10'sd7;
		12'd110: coeff = 10'sd8;
		12'd111: coeff = 10'sd8;
		12'd112: coeff = 10'sd8;
		12'd113: coeff = 10'sd8;
		12'd114: coeff = 10'sd8;
		12'd115: coeff = 10'sd8;
		12'd116: coeff = 10'sd8;
		12'd117: coeff = 10'sd9;
		12'd118: coeff = 10'sd9;
		12'd119: coeff = 10'sd9;
		12'd120: coeff = 10'sd9;
		12'd121: coeff = 10'sd9;
		12'd122: coeff = 10'sd9;
		12'd123: coeff = 10'sd10;
		12'd124: coeff = 10'sd10;
		12'd125: coeff = 10'sd10;
		12'd126: coeff = 10'sd10;
		12'd127: coeff = 10'sd10;
		12'd128: coeff = 10'sd10;
		12'd129: coeff = 10'sd10;
		12'd130: coeff = 10'sd11;
		12'd131: coeff = 10'sd11;
		12'd132: coeff = 10'sd11;
		12'd133: coeff = 10'sd11;
		12'd134: coeff = 10'sd11;
		12'd135: coeff = 10'sd11;
		12'd136: coeff = 10'sd12;
		12'd137: coeff = 10'sd12;
		12'd138: coeff = 10'sd12;
		12'd139: coeff = 10'sd12;
		12'd140: coeff = 10'sd12;
		12'd141: coeff = 10'sd13;
		12'd142: coeff = 10'sd13;
		12'd143: coeff = 10'sd13;
		12'd144: coeff = 10'sd13;
		12'd145: coeff = 10'sd13;
		12'd146: coeff = 10'sd13;
		12'd147: coeff = 10'sd14;
		12'd148: coeff = 10'sd14;
		12'd149: coeff = 10'sd14;
		12'd150: coeff = 10'sd14;
		12'd151: coeff = 10'sd14;
		12'd152: coeff = 10'sd15;
		12'd153: coeff = 10'sd15;
		12'd154: coeff = 10'sd15;
		12'd155: coeff = 10'sd15;
		12'd156: coeff = 10'sd15;
		12'd157: coeff = 10'sd15;
		12'd158: coeff = 10'sd16;
		12'd159: coeff = 10'sd16;
		12'd160: coeff = 10'sd16;
		12'd161: coeff = 10'sd16;
		12'd162: coeff = 10'sd16;
		12'd163: coeff = 10'sd17;
		12'd164: coeff = 10'sd17;
		12'd165: coeff = 10'sd17;
		12'd166: coeff = 10'sd17;
		12'd167: coeff = 10'sd18;
		12'd168: coeff = 10'sd18;
		12'd169: coeff = 10'sd18;
		12'd170: coeff = 10'sd18;
		12'd171: coeff = 10'sd18;
		12'd172: coeff = 10'sd19;
		12'd173: coeff = 10'sd19;
		12'd174: coeff = 10'sd19;
		12'd175: coeff = 10'sd19;
		12'd176: coeff = 10'sd19;
		12'd177: coeff = 10'sd20;
		12'd178: coeff = 10'sd20;
		12'd179: coeff = 10'sd20;
		12'd180: coeff = 10'sd20;
		12'd181: coeff = 10'sd21;
		12'd182: coeff = 10'sd21;
		12'd183: coeff = 10'sd21;
		12'd184: coeff = 10'sd21;
		12'd185: coeff = 10'sd21;
		12'd186: coeff = 10'sd22;
		12'd187: coeff = 10'sd22;
		12'd188: coeff = 10'sd22;
		12'd189: coeff = 10'sd22;
		12'd190: coeff = 10'sd23;
		12'd191: coeff = 10'sd23;
		12'd192: coeff = 10'sd23;
		12'd193: coeff = 10'sd23;
		12'd194: coeff = 10'sd24;
		12'd195: coeff = 10'sd24;
		12'd196: coeff = 10'sd24;
		12'd197: coeff = 10'sd24;
		12'd198: coeff = 10'sd25;
		12'd199: coeff = 10'sd25;
		12'd200: coeff = 10'sd25;
		12'd201: coeff = 10'sd25;
		12'd202: coeff = 10'sd26;
		12'd203: coeff = 10'sd26;
		12'd204: coeff = 10'sd26;
		12'd205: coeff = 10'sd26;
		12'd206: coeff = 10'sd27;
		12'd207: coeff = 10'sd27;
		12'd208: coeff = 10'sd27;
		12'd209: coeff = 10'sd27;
		12'd210: coeff = 10'sd28;
		12'd211: coeff = 10'sd28;
		12'd212: coeff = 10'sd28;
		12'd213: coeff = 10'sd28;
		12'd214: coeff = 10'sd29;
		12'd215: coeff = 10'sd29;
		12'd216: coeff = 10'sd29;
		12'd217: coeff = 10'sd29;
		12'd218: coeff = 10'sd30;
		12'd219: coeff = 10'sd30;
		12'd220: coeff = 10'sd30;
		12'd221: coeff = 10'sd31;
		12'd222: coeff = 10'sd31;
		12'd223: coeff = 10'sd31;
		12'd224: coeff = 10'sd31;
		12'd225: coeff = 10'sd32;
		12'd226: coeff = 10'sd32;
		12'd227: coeff = 10'sd32;
		12'd228: coeff = 10'sd33;
		12'd229: coeff = 10'sd33;
		12'd230: coeff = 10'sd33;
		12'd231: coeff = 10'sd33;
		12'd232: coeff = 10'sd34;
		12'd233: coeff = 10'sd34;
		12'd234: coeff = 10'sd34;
		12'd235: coeff = 10'sd35;
		12'd236: coeff = 10'sd35;
		12'd237: coeff = 10'sd35;
		12'd238: coeff = 10'sd35;
		12'd239: coeff = 10'sd36;
		12'd240: coeff = 10'sd36;
		12'd241: coeff = 10'sd36;
		12'd242: coeff = 10'sd37;
		12'd243: coeff = 10'sd37;
		12'd244: coeff = 10'sd37;
		12'd245: coeff = 10'sd37;
		12'd246: coeff = 10'sd38;
		12'd247: coeff = 10'sd38;
		12'd248: coeff = 10'sd38;
		12'd249: coeff = 10'sd39;
		12'd250: coeff = 10'sd39;
		12'd251: coeff = 10'sd39;
		12'd252: coeff = 10'sd40;
		12'd253: coeff = 10'sd40;
		12'd254: coeff = 10'sd40;
		12'd255: coeff = 10'sd41;
		12'd256: coeff = 10'sd41;
		12'd257: coeff = 10'sd41;
		12'd258: coeff = 10'sd41;
		12'd259: coeff = 10'sd42;
		12'd260: coeff = 10'sd42;
		12'd261: coeff = 10'sd42;
		12'd262: coeff = 10'sd43;
		12'd263: coeff = 10'sd43;
		12'd264: coeff = 10'sd43;
		12'd265: coeff = 10'sd44;
		12'd266: coeff = 10'sd44;
		12'd267: coeff = 10'sd44;
		12'd268: coeff = 10'sd45;
		12'd269: coeff = 10'sd45;
		12'd270: coeff = 10'sd45;
		12'd271: coeff = 10'sd46;
		12'd272: coeff = 10'sd46;
		12'd273: coeff = 10'sd46;
		12'd274: coeff = 10'sd47;
		12'd275: coeff = 10'sd47;
		12'd276: coeff = 10'sd47;
		12'd277: coeff = 10'sd48;
		12'd278: coeff = 10'sd48;
		12'd279: coeff = 10'sd48;
		12'd280: coeff = 10'sd49;
		12'd281: coeff = 10'sd49;
		12'd282: coeff = 10'sd49;
		12'd283: coeff = 10'sd50;
		12'd284: coeff = 10'sd50;
		12'd285: coeff = 10'sd50;
		12'd286: coeff = 10'sd51;
		12'd287: coeff = 10'sd51;
		12'd288: coeff = 10'sd52;
		12'd289: coeff = 10'sd52;
		12'd290: coeff = 10'sd52;
		12'd291: coeff = 10'sd53;
		12'd292: coeff = 10'sd53;
		12'd293: coeff = 10'sd53;
		12'd294: coeff = 10'sd54;
		12'd295: coeff = 10'sd54;
		12'd296: coeff = 10'sd54;
		12'd297: coeff = 10'sd55;
		12'd298: coeff = 10'sd55;
		12'd299: coeff = 10'sd55;
		12'd300: coeff = 10'sd56;
		12'd301: coeff = 10'sd56;
		12'd302: coeff = 10'sd57;
		12'd303: coeff = 10'sd57;
		12'd304: coeff = 10'sd57;
		12'd305: coeff = 10'sd58;
		12'd306: coeff = 10'sd58;
		12'd307: coeff = 10'sd58;
		12'd308: coeff = 10'sd59;
		12'd309: coeff = 10'sd59;
		12'd310: coeff = 10'sd60;
		12'd311: coeff = 10'sd60;
		12'd312: coeff = 10'sd60;
		12'd313: coeff = 10'sd61;
		12'd314: coeff = 10'sd61;
		12'd315: coeff = 10'sd61;
		12'd316: coeff = 10'sd62;
		12'd317: coeff = 10'sd62;
		12'd318: coeff = 10'sd63;
		12'd319: coeff = 10'sd63;
		12'd320: coeff = 10'sd63;
		12'd321: coeff = 10'sd64;
		12'd322: coeff = 10'sd64;
		12'd323: coeff = 10'sd65;
		12'd324: coeff = 10'sd65;
		12'd325: coeff = 10'sd65;
		12'd326: coeff = 10'sd66;
		12'd327: coeff = 10'sd66;
		12'd328: coeff = 10'sd66;
		12'd329: coeff = 10'sd67;
		12'd330: coeff = 10'sd67;
		12'd331: coeff = 10'sd68;
		12'd332: coeff = 10'sd68;
		12'd333: coeff = 10'sd68;
		12'd334: coeff = 10'sd69;
		12'd335: coeff = 10'sd69;
		12'd336: coeff = 10'sd70;
		12'd337: coeff = 10'sd70;
		12'd338: coeff = 10'sd71;
		12'd339: coeff = 10'sd71;
		12'd340: coeff = 10'sd71;
		12'd341: coeff = 10'sd72;
		12'd342: coeff = 10'sd72;
		12'd343: coeff = 10'sd73;
		12'd344: coeff = 10'sd73;
		12'd345: coeff = 10'sd73;
		12'd346: coeff = 10'sd74;
		12'd347: coeff = 10'sd74;
		12'd348: coeff = 10'sd75;
		12'd349: coeff = 10'sd75;
		12'd350: coeff = 10'sd75;
		12'd351: coeff = 10'sd76;
		12'd352: coeff = 10'sd76;
		12'd353: coeff = 10'sd77;
		12'd354: coeff = 10'sd77;
		12'd355: coeff = 10'sd78;
		12'd356: coeff = 10'sd78;
		12'd357: coeff = 10'sd78;
		12'd358: coeff = 10'sd79;
		12'd359: coeff = 10'sd79;
		12'd360: coeff = 10'sd80;
		12'd361: coeff = 10'sd80;
		12'd362: coeff = 10'sd81;
		12'd363: coeff = 10'sd81;
		12'd364: coeff = 10'sd81;
		12'd365: coeff = 10'sd82;
		12'd366: coeff = 10'sd82;
		12'd367: coeff = 10'sd83;
		12'd368: coeff = 10'sd83;
		12'd369: coeff = 10'sd84;
		12'd370: coeff = 10'sd84;
		12'd371: coeff = 10'sd85;
		12'd372: coeff = 10'sd85;
		12'd373: coeff = 10'sd85;
		12'd374: coeff = 10'sd86;
		12'd375: coeff = 10'sd86;
		12'd376: coeff = 10'sd87;
		12'd377: coeff = 10'sd87;
		12'd378: coeff = 10'sd88;
		12'd379: coeff = 10'sd88;
		12'd380: coeff = 10'sd89;
		12'd381: coeff = 10'sd89;
		12'd382: coeff = 10'sd89;
		12'd383: coeff = 10'sd90;
		12'd384: coeff = 10'sd90;
		12'd385: coeff = 10'sd91;
		12'd386: coeff = 10'sd91;
		12'd387: coeff = 10'sd92;
		12'd388: coeff = 10'sd92;
		12'd389: coeff = 10'sd93;
		12'd390: coeff = 10'sd93;
		12'd391: coeff = 10'sd94;
		12'd392: coeff = 10'sd94;
		12'd393: coeff = 10'sd95;
		12'd394: coeff = 10'sd95;
		12'd395: coeff = 10'sd95;
		12'd396: coeff = 10'sd96;
		12'd397: coeff = 10'sd96;
		12'd398: coeff = 10'sd97;
		12'd399: coeff = 10'sd97;
		12'd400: coeff = 10'sd98;
		12'd401: coeff = 10'sd98;
		12'd402: coeff = 10'sd99;
		12'd403: coeff = 10'sd99;
		12'd404: coeff = 10'sd100;
		12'd405: coeff = 10'sd100;
		12'd406: coeff = 10'sd101;
		12'd407: coeff = 10'sd101;
		12'd408: coeff = 10'sd102;
		12'd409: coeff = 10'sd102;
		12'd410: coeff = 10'sd103;
		12'd411: coeff = 10'sd103;
		12'd412: coeff = 10'sd104;
		12'd413: coeff = 10'sd104;
		12'd414: coeff = 10'sd105;
		12'd415: coeff = 10'sd105;
		12'd416: coeff = 10'sd106;
		12'd417: coeff = 10'sd106;
		12'd418: coeff = 10'sd107;
		12'd419: coeff = 10'sd107;
		12'd420: coeff = 10'sd107;
		12'd421: coeff = 10'sd108;
		12'd422: coeff = 10'sd108;
		12'd423: coeff = 10'sd109;
		12'd424: coeff = 10'sd109;
		12'd425: coeff = 10'sd110;
		12'd426: coeff = 10'sd110;
		12'd427: coeff = 10'sd111;
		12'd428: coeff = 10'sd111;
		12'd429: coeff = 10'sd112;
		12'd430: coeff = 10'sd112;
		12'd431: coeff = 10'sd113;
		12'd432: coeff = 10'sd113;
		12'd433: coeff = 10'sd114;
		12'd434: coeff = 10'sd114;
		12'd435: coeff = 10'sd115;
		12'd436: coeff = 10'sd116;
		12'd437: coeff = 10'sd116;
		12'd438: coeff = 10'sd117;
		12'd439: coeff = 10'sd117;
		12'd440: coeff = 10'sd118;
		12'd441: coeff = 10'sd118;
		12'd442: coeff = 10'sd119;
		12'd443: coeff = 10'sd119;
		12'd444: coeff = 10'sd120;
		12'd445: coeff = 10'sd120;
		12'd446: coeff = 10'sd121;
		12'd447: coeff = 10'sd121;
		12'd448: coeff = 10'sd122;
		12'd449: coeff = 10'sd122;
		12'd450: coeff = 10'sd123;
		12'd451: coeff = 10'sd123;
		12'd452: coeff = 10'sd124;
		12'd453: coeff = 10'sd124;
		12'd454: coeff = 10'sd125;
		12'd455: coeff = 10'sd125;
		12'd456: coeff = 10'sd126;
		12'd457: coeff = 10'sd126;
		12'd458: coeff = 10'sd127;
		12'd459: coeff = 10'sd127;
		12'd460: coeff = 10'sd128;
		12'd461: coeff = 10'sd129;
		12'd462: coeff = 10'sd129;
		12'd463: coeff = 10'sd130;
		12'd464: coeff = 10'sd130;
		12'd465: coeff = 10'sd131;
		12'd466: coeff = 10'sd131;
		12'd467: coeff = 10'sd132;
		12'd468: coeff = 10'sd132;
		12'd469: coeff = 10'sd133;
		12'd470: coeff = 10'sd133;
		12'd471: coeff = 10'sd134;
		12'd472: coeff = 10'sd134;
		12'd473: coeff = 10'sd135;
		12'd474: coeff = 10'sd136;
		12'd475: coeff = 10'sd136;
		12'd476: coeff = 10'sd137;
		12'd477: coeff = 10'sd137;
		12'd478: coeff = 10'sd138;
		12'd479: coeff = 10'sd138;
		12'd480: coeff = 10'sd139;
		12'd481: coeff = 10'sd139;
		12'd482: coeff = 10'sd140;
		12'd483: coeff = 10'sd140;
		12'd484: coeff = 10'sd141;
		12'd485: coeff = 10'sd142;
		12'd486: coeff = 10'sd142;
		12'd487: coeff = 10'sd143;
		12'd488: coeff = 10'sd143;
		12'd489: coeff = 10'sd144;
		12'd490: coeff = 10'sd144;
		12'd491: coeff = 10'sd145;
		12'd492: coeff = 10'sd146;
		12'd493: coeff = 10'sd146;
		12'd494: coeff = 10'sd147;
		12'd495: coeff = 10'sd147;
		12'd496: coeff = 10'sd148;
		12'd497: coeff = 10'sd148;
		12'd498: coeff = 10'sd149;
		12'd499: coeff = 10'sd149;
		12'd500: coeff = 10'sd150;
		12'd501: coeff = 10'sd151;
		12'd502: coeff = 10'sd151;
		12'd503: coeff = 10'sd152;
		12'd504: coeff = 10'sd152;
		12'd505: coeff = 10'sd153;
		12'd506: coeff = 10'sd153;
		12'd507: coeff = 10'sd154;
		12'd508: coeff = 10'sd155;
		12'd509: coeff = 10'sd155;
		12'd510: coeff = 10'sd156;
		12'd511: coeff = 10'sd156;
		12'd512: coeff = 10'sd157;
		12'd513: coeff = 10'sd158;
		12'd514: coeff = 10'sd158;
		12'd515: coeff = 10'sd159;
		12'd516: coeff = 10'sd159;
		12'd517: coeff = 10'sd160;
		12'd518: coeff = 10'sd160;
		12'd519: coeff = 10'sd161;
		12'd520: coeff = 10'sd162;
		12'd521: coeff = 10'sd162;
		12'd522: coeff = 10'sd163;
		12'd523: coeff = 10'sd163;
		12'd524: coeff = 10'sd164;
		12'd525: coeff = 10'sd165;
		12'd526: coeff = 10'sd165;
		12'd527: coeff = 10'sd166;
		12'd528: coeff = 10'sd166;
		12'd529: coeff = 10'sd167;
		12'd530: coeff = 10'sd167;
		12'd531: coeff = 10'sd168;
		12'd532: coeff = 10'sd169;
		12'd533: coeff = 10'sd169;
		12'd534: coeff = 10'sd170;
		12'd535: coeff = 10'sd170;
		12'd536: coeff = 10'sd171;
		12'd537: coeff = 10'sd172;
		12'd538: coeff = 10'sd172;
		12'd539: coeff = 10'sd173;
		12'd540: coeff = 10'sd173;
		12'd541: coeff = 10'sd174;
		12'd542: coeff = 10'sd175;
		12'd543: coeff = 10'sd175;
		12'd544: coeff = 10'sd176;
		12'd545: coeff = 10'sd177;
		12'd546: coeff = 10'sd177;
		12'd547: coeff = 10'sd178;
		12'd548: coeff = 10'sd178;
		12'd549: coeff = 10'sd179;
		12'd550: coeff = 10'sd180;
		12'd551: coeff = 10'sd180;
		12'd552: coeff = 10'sd181;
		12'd553: coeff = 10'sd181;
		12'd554: coeff = 10'sd182;
		12'd555: coeff = 10'sd183;
		12'd556: coeff = 10'sd183;
		12'd557: coeff = 10'sd184;
		12'd558: coeff = 10'sd184;
		12'd559: coeff = 10'sd185;
		12'd560: coeff = 10'sd186;
		12'd561: coeff = 10'sd186;
		12'd562: coeff = 10'sd187;
		12'd563: coeff = 10'sd188;
		12'd564: coeff = 10'sd188;
		12'd565: coeff = 10'sd189;
		12'd566: coeff = 10'sd189;
		12'd567: coeff = 10'sd190;
		12'd568: coeff = 10'sd191;
		12'd569: coeff = 10'sd191;
		12'd570: coeff = 10'sd192;
		12'd571: coeff = 10'sd193;
		12'd572: coeff = 10'sd193;
		12'd573: coeff = 10'sd194;
		12'd574: coeff = 10'sd194;
		12'd575: coeff = 10'sd195;
		12'd576: coeff = 10'sd196;
		12'd577: coeff = 10'sd196;
		12'd578: coeff = 10'sd197;
		12'd579: coeff = 10'sd198;
		12'd580: coeff = 10'sd198;
		12'd581: coeff = 10'sd199;
		12'd582: coeff = 10'sd200;
		12'd583: coeff = 10'sd200;
		12'd584: coeff = 10'sd201;
		12'd585: coeff = 10'sd201;
		12'd586: coeff = 10'sd202;
		12'd587: coeff = 10'sd203;
		12'd588: coeff = 10'sd203;
		12'd589: coeff = 10'sd204;
		12'd590: coeff = 10'sd205;
		12'd591: coeff = 10'sd205;
		12'd592: coeff = 10'sd206;
		12'd593: coeff = 10'sd207;
		12'd594: coeff = 10'sd207;
		12'd595: coeff = 10'sd208;
		12'd596: coeff = 10'sd209;
		12'd597: coeff = 10'sd209;
		12'd598: coeff = 10'sd210;
		12'd599: coeff = 10'sd211;
		12'd600: coeff = 10'sd211;
		12'd601: coeff = 10'sd212;
		12'd602: coeff = 10'sd212;
		12'd603: coeff = 10'sd213;
		12'd604: coeff = 10'sd214;
		12'd605: coeff = 10'sd214;
		12'd606: coeff = 10'sd215;
		12'd607: coeff = 10'sd216;
		12'd608: coeff = 10'sd216;
		12'd609: coeff = 10'sd217;
		12'd610: coeff = 10'sd218;
		12'd611: coeff = 10'sd218;
		12'd612: coeff = 10'sd219;
		12'd613: coeff = 10'sd220;
		12'd614: coeff = 10'sd220;
		12'd615: coeff = 10'sd221;
		12'd616: coeff = 10'sd222;
		12'd617: coeff = 10'sd222;
		12'd618: coeff = 10'sd223;
		12'd619: coeff = 10'sd224;
		12'd620: coeff = 10'sd224;
		12'd621: coeff = 10'sd225;
		12'd622: coeff = 10'sd226;
		12'd623: coeff = 10'sd226;
		12'd624: coeff = 10'sd227;
		12'd625: coeff = 10'sd228;
		12'd626: coeff = 10'sd228;
		12'd627: coeff = 10'sd229;
		12'd628: coeff = 10'sd230;
		12'd629: coeff = 10'sd230;
		12'd630: coeff = 10'sd231;
		12'd631: coeff = 10'sd232;
		12'd632: coeff = 10'sd232;
		12'd633: coeff = 10'sd233;
		12'd634: coeff = 10'sd234;
		12'd635: coeff = 10'sd234;
		12'd636: coeff = 10'sd235;
		12'd637: coeff = 10'sd236;
		12'd638: coeff = 10'sd236;
		12'd639: coeff = 10'sd237;
		12'd640: coeff = 10'sd238;
		12'd641: coeff = 10'sd238;
		12'd642: coeff = 10'sd239;
		12'd643: coeff = 10'sd240;
		12'd644: coeff = 10'sd240;
		12'd645: coeff = 10'sd241;
		12'd646: coeff = 10'sd242;
		12'd647: coeff = 10'sd243;
		12'd648: coeff = 10'sd243;
		12'd649: coeff = 10'sd244;
		12'd650: coeff = 10'sd245;
		12'd651: coeff = 10'sd245;
		12'd652: coeff = 10'sd246;
		12'd653: coeff = 10'sd247;
		12'd654: coeff = 10'sd247;
		12'd655: coeff = 10'sd248;
		12'd656: coeff = 10'sd249;
		12'd657: coeff = 10'sd249;
		12'd658: coeff = 10'sd250;
		12'd659: coeff = 10'sd251;
		12'd660: coeff = 10'sd251;
		12'd661: coeff = 10'sd252;
		12'd662: coeff = 10'sd253;
		12'd663: coeff = 10'sd254;
		12'd664: coeff = 10'sd254;
		12'd665: coeff = 10'sd255;
		12'd666: coeff = 10'sd256;
		12'd667: coeff = 10'sd256;
		12'd668: coeff = 10'sd257;
		12'd669: coeff = 10'sd258;
		12'd670: coeff = 10'sd258;
		12'd671: coeff = 10'sd259;
		12'd672: coeff = 10'sd260;
		12'd673: coeff = 10'sd261;
		12'd674: coeff = 10'sd261;
		12'd675: coeff = 10'sd262;
		12'd676: coeff = 10'sd263;
		12'd677: coeff = 10'sd263;
		12'd678: coeff = 10'sd264;
		12'd679: coeff = 10'sd265;
		12'd680: coeff = 10'sd265;
		12'd681: coeff = 10'sd266;
		12'd682: coeff = 10'sd267;
		12'd683: coeff = 10'sd268;
		12'd684: coeff = 10'sd268;
		12'd685: coeff = 10'sd269;
		12'd686: coeff = 10'sd270;
		12'd687: coeff = 10'sd270;
		12'd688: coeff = 10'sd271;
		12'd689: coeff = 10'sd272;
		12'd690: coeff = 10'sd273;
		12'd691: coeff = 10'sd273;
		12'd692: coeff = 10'sd274;
		12'd693: coeff = 10'sd275;
		12'd694: coeff = 10'sd275;
		12'd695: coeff = 10'sd276;
		12'd696: coeff = 10'sd277;
		12'd697: coeff = 10'sd278;
		12'd698: coeff = 10'sd278;
		12'd699: coeff = 10'sd279;
		12'd700: coeff = 10'sd280;
		12'd701: coeff = 10'sd280;
		12'd702: coeff = 10'sd281;
		12'd703: coeff = 10'sd282;
		12'd704: coeff = 10'sd283;
		12'd705: coeff = 10'sd283;
		12'd706: coeff = 10'sd284;
		12'd707: coeff = 10'sd285;
		12'd708: coeff = 10'sd285;
		12'd709: coeff = 10'sd286;
		12'd710: coeff = 10'sd287;
		12'd711: coeff = 10'sd288;
		12'd712: coeff = 10'sd288;
		12'd713: coeff = 10'sd289;
		12'd714: coeff = 10'sd290;
		12'd715: coeff = 10'sd290;
		12'd716: coeff = 10'sd291;
		12'd717: coeff = 10'sd292;
		12'd718: coeff = 10'sd293;
		12'd719: coeff = 10'sd293;
		12'd720: coeff = 10'sd294;
		12'd721: coeff = 10'sd295;
		12'd722: coeff = 10'sd296;
		12'd723: coeff = 10'sd296;
		12'd724: coeff = 10'sd297;
		12'd725: coeff = 10'sd298;
		12'd726: coeff = 10'sd299;
		12'd727: coeff = 10'sd299;
		12'd728: coeff = 10'sd300;
		12'd729: coeff = 10'sd301;
		12'd730: coeff = 10'sd301;
		12'd731: coeff = 10'sd302;
		12'd732: coeff = 10'sd303;
		12'd733: coeff = 10'sd304;
		12'd734: coeff = 10'sd304;
		12'd735: coeff = 10'sd305;
		12'd736: coeff = 10'sd306;
		12'd737: coeff = 10'sd307;
		12'd738: coeff = 10'sd307;
		12'd739: coeff = 10'sd308;
		12'd740: coeff = 10'sd309;
		12'd741: coeff = 10'sd310;
		12'd742: coeff = 10'sd310;
		12'd743: coeff = 10'sd311;
		12'd744: coeff = 10'sd312;
		12'd745: coeff = 10'sd312;
		12'd746: coeff = 10'sd313;
		12'd747: coeff = 10'sd314;
		12'd748: coeff = 10'sd315;
		12'd749: coeff = 10'sd315;
		12'd750: coeff = 10'sd316;
		12'd751: coeff = 10'sd317;
		12'd752: coeff = 10'sd318;
		12'd753: coeff = 10'sd318;
		12'd754: coeff = 10'sd319;
		12'd755: coeff = 10'sd320;
		12'd756: coeff = 10'sd321;
		12'd757: coeff = 10'sd321;
		12'd758: coeff = 10'sd322;
		12'd759: coeff = 10'sd323;
		12'd760: coeff = 10'sd324;
		12'd761: coeff = 10'sd324;
		12'd762: coeff = 10'sd325;
		12'd763: coeff = 10'sd326;
		12'd764: coeff = 10'sd327;
		12'd765: coeff = 10'sd327;
		12'd766: coeff = 10'sd328;
		12'd767: coeff = 10'sd329;
		12'd768: coeff = 10'sd330;
		12'd769: coeff = 10'sd330;
		12'd770: coeff = 10'sd331;
		12'd771: coeff = 10'sd332;
		12'd772: coeff = 10'sd333;
		12'd773: coeff = 10'sd333;
		12'd774: coeff = 10'sd334;
		12'd775: coeff = 10'sd335;
		12'd776: coeff = 10'sd336;
		12'd777: coeff = 10'sd336;
		12'd778: coeff = 10'sd337;
		12'd779: coeff = 10'sd338;
		12'd780: coeff = 10'sd339;
		12'd781: coeff = 10'sd339;
		12'd782: coeff = 10'sd340;
		12'd783: coeff = 10'sd341;
		12'd784: coeff = 10'sd342;
		12'd785: coeff = 10'sd343;
		12'd786: coeff = 10'sd343;
		12'd787: coeff = 10'sd344;
		12'd788: coeff = 10'sd345;
		12'd789: coeff = 10'sd346;
		12'd790: coeff = 10'sd346;
		12'd791: coeff = 10'sd347;
		12'd792: coeff = 10'sd348;
		12'd793: coeff = 10'sd349;
		12'd794: coeff = 10'sd349;
		12'd795: coeff = 10'sd350;
		12'd796: coeff = 10'sd351;
		12'd797: coeff = 10'sd352;
		12'd798: coeff = 10'sd352;
		12'd799: coeff = 10'sd353;
		12'd800: coeff = 10'sd354;
		12'd801: coeff = 10'sd355;
		12'd802: coeff = 10'sd355;
		12'd803: coeff = 10'sd356;
		12'd804: coeff = 10'sd357;
		12'd805: coeff = 10'sd358;
		12'd806: coeff = 10'sd359;
		12'd807: coeff = 10'sd359;
		12'd808: coeff = 10'sd360;
		12'd809: coeff = 10'sd361;
		12'd810: coeff = 10'sd362;
		12'd811: coeff = 10'sd362;
		12'd812: coeff = 10'sd363;
		12'd813: coeff = 10'sd364;
		12'd814: coeff = 10'sd365;
		12'd815: coeff = 10'sd365;
		12'd816: coeff = 10'sd366;
		12'd817: coeff = 10'sd367;
		12'd818: coeff = 10'sd368;
		12'd819: coeff = 10'sd369;
		12'd820: coeff = 10'sd369;
		12'd821: coeff = 10'sd370;
		12'd822: coeff = 10'sd371;
		12'd823: coeff = 10'sd372;
		12'd824: coeff = 10'sd372;
		12'd825: coeff = 10'sd373;
		12'd826: coeff = 10'sd374;
		12'd827: coeff = 10'sd375;
		12'd828: coeff = 10'sd376;
		12'd829: coeff = 10'sd376;
		12'd830: coeff = 10'sd377;
		12'd831: coeff = 10'sd378;
		12'd832: coeff = 10'sd379;
		12'd833: coeff = 10'sd379;
		12'd834: coeff = 10'sd380;
		12'd835: coeff = 10'sd381;
		12'd836: coeff = 10'sd382;
		12'd837: coeff = 10'sd382;
		12'd838: coeff = 10'sd383;
		12'd839: coeff = 10'sd384;
		12'd840: coeff = 10'sd385;
		12'd841: coeff = 10'sd386;
		12'd842: coeff = 10'sd386;
		12'd843: coeff = 10'sd387;
		12'd844: coeff = 10'sd388;
		12'd845: coeff = 10'sd389;
		12'd846: coeff = 10'sd390;
		12'd847: coeff = 10'sd390;
		12'd848: coeff = 10'sd391;
		12'd849: coeff = 10'sd392;
		12'd850: coeff = 10'sd393;
		12'd851: coeff = 10'sd393;
		12'd852: coeff = 10'sd394;
		12'd853: coeff = 10'sd395;
		12'd854: coeff = 10'sd396;
		12'd855: coeff = 10'sd397;
		12'd856: coeff = 10'sd397;
		12'd857: coeff = 10'sd398;
		12'd858: coeff = 10'sd399;
		12'd859: coeff = 10'sd400;
		12'd860: coeff = 10'sd400;
		12'd861: coeff = 10'sd401;
		12'd862: coeff = 10'sd402;
		12'd863: coeff = 10'sd403;
		12'd864: coeff = 10'sd404;
		12'd865: coeff = 10'sd404;
		12'd866: coeff = 10'sd405;
		12'd867: coeff = 10'sd406;
		12'd868: coeff = 10'sd407;
		12'd869: coeff = 10'sd408;
		12'd870: coeff = 10'sd408;
		12'd871: coeff = 10'sd409;
		12'd872: coeff = 10'sd410;
		12'd873: coeff = 10'sd411;
		12'd874: coeff = 10'sd411;
		12'd875: coeff = 10'sd412;
		12'd876: coeff = 10'sd413;
		12'd877: coeff = 10'sd414;
		12'd878: coeff = 10'sd415;
		12'd879: coeff = 10'sd415;
		12'd880: coeff = 10'sd416;
		12'd881: coeff = 10'sd417;
		12'd882: coeff = 10'sd418;
		12'd883: coeff = 10'sd419;
		12'd884: coeff = 10'sd419;
		12'd885: coeff = 10'sd420;
		12'd886: coeff = 10'sd421;
		12'd887: coeff = 10'sd422;
		12'd888: coeff = 10'sd423;
		12'd889: coeff = 10'sd423;
		12'd890: coeff = 10'sd424;
		12'd891: coeff = 10'sd425;
		12'd892: coeff = 10'sd426;
		12'd893: coeff = 10'sd427;
		12'd894: coeff = 10'sd427;
		12'd895: coeff = 10'sd428;
		12'd896: coeff = 10'sd429;
		12'd897: coeff = 10'sd430;
		12'd898: coeff = 10'sd430;
		12'd899: coeff = 10'sd431;
		12'd900: coeff = 10'sd432;
		12'd901: coeff = 10'sd433;
		12'd902: coeff = 10'sd434;
		12'd903: coeff = 10'sd434;
		12'd904: coeff = 10'sd435;
		12'd905: coeff = 10'sd436;
		12'd906: coeff = 10'sd437;
		12'd907: coeff = 10'sd438;
		12'd908: coeff = 10'sd438;
		12'd909: coeff = 10'sd439;
		12'd910: coeff = 10'sd440;
		12'd911: coeff = 10'sd441;
		12'd912: coeff = 10'sd442;
		12'd913: coeff = 10'sd442;
		12'd914: coeff = 10'sd443;
		12'd915: coeff = 10'sd444;
		12'd916: coeff = 10'sd445;
		12'd917: coeff = 10'sd446;
		12'd918: coeff = 10'sd446;
		12'd919: coeff = 10'sd447;
		12'd920: coeff = 10'sd448;
		12'd921: coeff = 10'sd449;
		12'd922: coeff = 10'sd450;
		12'd923: coeff = 10'sd450;
		12'd924: coeff = 10'sd451;
		12'd925: coeff = 10'sd452;
		12'd926: coeff = 10'sd453;
		12'd927: coeff = 10'sd454;
		12'd928: coeff = 10'sd454;
		12'd929: coeff = 10'sd455;
		12'd930: coeff = 10'sd456;
		12'd931: coeff = 10'sd457;
		12'd932: coeff = 10'sd458;
		12'd933: coeff = 10'sd458;
		12'd934: coeff = 10'sd459;
		12'd935: coeff = 10'sd460;
		12'd936: coeff = 10'sd461;
		12'd937: coeff = 10'sd462;
		12'd938: coeff = 10'sd462;
		12'd939: coeff = 10'sd463;
		12'd940: coeff = 10'sd464;
		12'd941: coeff = 10'sd465;
		12'd942: coeff = 10'sd466;
		12'd943: coeff = 10'sd466;
		12'd944: coeff = 10'sd467;
		12'd945: coeff = 10'sd468;
		12'd946: coeff = 10'sd469;
		12'd947: coeff = 10'sd470;
		12'd948: coeff = 10'sd470;
		12'd949: coeff = 10'sd471;
		12'd950: coeff = 10'sd472;
		12'd951: coeff = 10'sd473;
		12'd952: coeff = 10'sd474;
		12'd953: coeff = 10'sd474;
		12'd954: coeff = 10'sd475;
		12'd955: coeff = 10'sd476;
		12'd956: coeff = 10'sd477;
		12'd957: coeff = 10'sd478;
		12'd958: coeff = 10'sd478;
		12'd959: coeff = 10'sd479;
		12'd960: coeff = 10'sd480;
		12'd961: coeff = 10'sd481;
		12'd962: coeff = 10'sd482;
		12'd963: coeff = 10'sd482;
		12'd964: coeff = 10'sd483;
		12'd965: coeff = 10'sd484;
		12'd966: coeff = 10'sd485;
		12'd967: coeff = 10'sd486;
		12'd968: coeff = 10'sd486;
		12'd969: coeff = 10'sd487;
		12'd970: coeff = 10'sd488;
		12'd971: coeff = 10'sd489;
		12'd972: coeff = 10'sd490;
		12'd973: coeff = 10'sd490;
		12'd974: coeff = 10'sd491;
		12'd975: coeff = 10'sd492;
		12'd976: coeff = 10'sd493;
		12'd977: coeff = 10'sd494;
		12'd978: coeff = 10'sd495;
		12'd979: coeff = 10'sd495;
		12'd980: coeff = 10'sd496;
		12'd981: coeff = 10'sd497;
		12'd982: coeff = 10'sd498;
		12'd983: coeff = 10'sd499;
		12'd984: coeff = 10'sd499;
		12'd985: coeff = 10'sd500;
		12'd986: coeff = 10'sd501;
		12'd987: coeff = 10'sd502;
		12'd988: coeff = 10'sd503;
		12'd989: coeff = 10'sd503;
		12'd990: coeff = 10'sd504;
		12'd991: coeff = 10'sd505;
		12'd992: coeff = 10'sd506;
		12'd993: coeff = 10'sd507;
		12'd994: coeff = 10'sd507;
		12'd995: coeff = 10'sd508;
		12'd996: coeff = 10'sd509;
		12'd997: coeff = 10'sd510;
		12'd998: coeff = 10'sd511;
		12'd999: coeff = 10'sd511;
		12'd1000: coeff = 10'sd512;
		12'd1001: coeff = 10'sd513;
		12'd1002: coeff = 10'sd514;
		12'd1003: coeff = 10'sd515;
		12'd1004: coeff = 10'sd515;
		12'd1005: coeff = 10'sd516;
		12'd1006: coeff = 10'sd517;
		12'd1007: coeff = 10'sd518;
		12'd1008: coeff = 10'sd519;
		12'd1009: coeff = 10'sd519;
		12'd1010: coeff = 10'sd520;
		12'd1011: coeff = 10'sd521;
		12'd1012: coeff = 10'sd522;
		12'd1013: coeff = 10'sd523;
		12'd1014: coeff = 10'sd523;
		12'd1015: coeff = 10'sd524;
		12'd1016: coeff = 10'sd525;
		12'd1017: coeff = 10'sd526;
		12'd1018: coeff = 10'sd527;
		12'd1019: coeff = 10'sd527;
		12'd1020: coeff = 10'sd528;
		12'd1021: coeff = 10'sd529;
		12'd1022: coeff = 10'sd530;
		12'd1023: coeff = 10'sd531;
		12'd1024: coeff = 10'sd532;
		12'd1025: coeff = 10'sd532;
		12'd1026: coeff = 10'sd533;
		12'd1027: coeff = 10'sd534;
		12'd1028: coeff = 10'sd535;
		12'd1029: coeff = 10'sd536;
		12'd1030: coeff = 10'sd536;
		12'd1031: coeff = 10'sd537;
		12'd1032: coeff = 10'sd538;
		12'd1033: coeff = 10'sd539;
		12'd1034: coeff = 10'sd540;
		12'd1035: coeff = 10'sd540;
		12'd1036: coeff = 10'sd541;
		12'd1037: coeff = 10'sd542;
		12'd1038: coeff = 10'sd543;
		12'd1039: coeff = 10'sd544;
		12'd1040: coeff = 10'sd544;
		12'd1041: coeff = 10'sd545;
		12'd1042: coeff = 10'sd546;
		12'd1043: coeff = 10'sd547;
		12'd1044: coeff = 10'sd548;
		12'd1045: coeff = 10'sd548;
		12'd1046: coeff = 10'sd549;
		12'd1047: coeff = 10'sd550;
		12'd1048: coeff = 10'sd551;
		12'd1049: coeff = 10'sd552;
		12'd1050: coeff = 10'sd552;
		12'd1051: coeff = 10'sd553;
		12'd1052: coeff = 10'sd554;
		12'd1053: coeff = 10'sd555;
		12'd1054: coeff = 10'sd556;
		12'd1055: coeff = 10'sd556;
		12'd1056: coeff = 10'sd557;
		12'd1057: coeff = 10'sd558;
		12'd1058: coeff = 10'sd559;
		12'd1059: coeff = 10'sd560;
		12'd1060: coeff = 10'sd560;
		12'd1061: coeff = 10'sd561;
		12'd1062: coeff = 10'sd562;
		12'd1063: coeff = 10'sd563;
		12'd1064: coeff = 10'sd564;
		12'd1065: coeff = 10'sd564;
		12'd1066: coeff = 10'sd565;
		12'd1067: coeff = 10'sd566;
		12'd1068: coeff = 10'sd567;
		12'd1069: coeff = 10'sd568;
		12'd1070: coeff = 10'sd568;
		12'd1071: coeff = 10'sd569;
		12'd1072: coeff = 10'sd570;
		12'd1073: coeff = 10'sd571;
		12'd1074: coeff = 10'sd572;
		12'd1075: coeff = 10'sd572;
		12'd1076: coeff = 10'sd573;
		12'd1077: coeff = 10'sd574;
		12'd1078: coeff = 10'sd575;
		12'd1079: coeff = 10'sd576;
		12'd1080: coeff = 10'sd576;
		12'd1081: coeff = 10'sd577;
		12'd1082: coeff = 10'sd578;
		12'd1083: coeff = 10'sd579;
		12'd1084: coeff = 10'sd580;
		12'd1085: coeff = 10'sd580;
		12'd1086: coeff = 10'sd581;
		12'd1087: coeff = 10'sd582;
		12'd1088: coeff = 10'sd583;
		12'd1089: coeff = 10'sd584;
		12'd1090: coeff = 10'sd584;
		12'd1091: coeff = 10'sd585;
		12'd1092: coeff = 10'sd586;
		12'd1093: coeff = 10'sd587;
		12'd1094: coeff = 10'sd588;
		12'd1095: coeff = 10'sd588;
		12'd1096: coeff = 10'sd589;
		12'd1097: coeff = 10'sd590;
		12'd1098: coeff = 10'sd591;
		12'd1099: coeff = 10'sd592;
		12'd1100: coeff = 10'sd592;
		12'd1101: coeff = 10'sd593;
		12'd1102: coeff = 10'sd594;
		12'd1103: coeff = 10'sd595;
		12'd1104: coeff = 10'sd595;
		12'd1105: coeff = 10'sd596;
		12'd1106: coeff = 10'sd597;
		12'd1107: coeff = 10'sd598;
		12'd1108: coeff = 10'sd599;
		12'd1109: coeff = 10'sd599;
		12'd1110: coeff = 10'sd600;
		12'd1111: coeff = 10'sd601;
		12'd1112: coeff = 10'sd602;
		12'd1113: coeff = 10'sd603;
		12'd1114: coeff = 10'sd603;
		12'd1115: coeff = 10'sd604;
		12'd1116: coeff = 10'sd605;
		12'd1117: coeff = 10'sd606;
		12'd1118: coeff = 10'sd607;
		12'd1119: coeff = 10'sd607;
		12'd1120: coeff = 10'sd608;
		12'd1121: coeff = 10'sd609;
		12'd1122: coeff = 10'sd610;
		12'd1123: coeff = 10'sd611;
		12'd1124: coeff = 10'sd611;
		12'd1125: coeff = 10'sd612;
		12'd1126: coeff = 10'sd613;
		12'd1127: coeff = 10'sd614;
		12'd1128: coeff = 10'sd614;
		12'd1129: coeff = 10'sd615;
		12'd1130: coeff = 10'sd616;
		12'd1131: coeff = 10'sd617;
		12'd1132: coeff = 10'sd618;
		12'd1133: coeff = 10'sd618;
		12'd1134: coeff = 10'sd619;
		12'd1135: coeff = 10'sd620;
		12'd1136: coeff = 10'sd621;
		12'd1137: coeff = 10'sd622;
		12'd1138: coeff = 10'sd622;
		12'd1139: coeff = 10'sd623;
		12'd1140: coeff = 10'sd624;
		12'd1141: coeff = 10'sd625;
		12'd1142: coeff = 10'sd625;
		12'd1143: coeff = 10'sd626;
		12'd1144: coeff = 10'sd627;
		12'd1145: coeff = 10'sd628;
		12'd1146: coeff = 10'sd629;
		12'd1147: coeff = 10'sd629;
		12'd1148: coeff = 10'sd630;
		12'd1149: coeff = 10'sd631;
		12'd1150: coeff = 10'sd632;
		12'd1151: coeff = 10'sd633;
		12'd1152: coeff = 10'sd633;
		12'd1153: coeff = 10'sd634;
		12'd1154: coeff = 10'sd635;
		12'd1155: coeff = 10'sd636;
		12'd1156: coeff = 10'sd636;
		12'd1157: coeff = 10'sd637;
		12'd1158: coeff = 10'sd638;
		12'd1159: coeff = 10'sd639;
		12'd1160: coeff = 10'sd640;
		12'd1161: coeff = 10'sd640;
		12'd1162: coeff = 10'sd641;
		12'd1163: coeff = 10'sd642;
		12'd1164: coeff = 10'sd643;
		12'd1165: coeff = 10'sd643;
		12'd1166: coeff = 10'sd644;
		12'd1167: coeff = 10'sd645;
		12'd1168: coeff = 10'sd646;
		12'd1169: coeff = 10'sd647;
		12'd1170: coeff = 10'sd647;
		12'd1171: coeff = 10'sd648;
		12'd1172: coeff = 10'sd649;
		12'd1173: coeff = 10'sd650;
		12'd1174: coeff = 10'sd650;
		12'd1175: coeff = 10'sd651;
		12'd1176: coeff = 10'sd652;
		12'd1177: coeff = 10'sd653;
		12'd1178: coeff = 10'sd654;
		12'd1179: coeff = 10'sd654;
		12'd1180: coeff = 10'sd655;
		12'd1181: coeff = 10'sd656;
		12'd1182: coeff = 10'sd657;
		12'd1183: coeff = 10'sd657;
		12'd1184: coeff = 10'sd658;
		12'd1185: coeff = 10'sd659;
		12'd1186: coeff = 10'sd660;
		12'd1187: coeff = 10'sd660;
		12'd1188: coeff = 10'sd661;
		12'd1189: coeff = 10'sd662;
		12'd1190: coeff = 10'sd663;
		12'd1191: coeff = 10'sd664;
		12'd1192: coeff = 10'sd664;
		12'd1193: coeff = 10'sd665;
		12'd1194: coeff = 10'sd666;
		12'd1195: coeff = 10'sd667;
		12'd1196: coeff = 10'sd667;
		12'd1197: coeff = 10'sd668;
		12'd1198: coeff = 10'sd669;
		12'd1199: coeff = 10'sd670;
		12'd1200: coeff = 10'sd670;
		12'd1201: coeff = 10'sd671;
		12'd1202: coeff = 10'sd672;
		12'd1203: coeff = 10'sd673;
		12'd1204: coeff = 10'sd674;
		12'd1205: coeff = 10'sd674;
		12'd1206: coeff = 10'sd675;
		12'd1207: coeff = 10'sd676;
		12'd1208: coeff = 10'sd677;
		12'd1209: coeff = 10'sd677;
		12'd1210: coeff = 10'sd678;
		12'd1211: coeff = 10'sd679;
		12'd1212: coeff = 10'sd680;
		12'd1213: coeff = 10'sd680;
		12'd1214: coeff = 10'sd681;
		12'd1215: coeff = 10'sd682;
		12'd1216: coeff = 10'sd683;
		12'd1217: coeff = 10'sd683;
		12'd1218: coeff = 10'sd684;
		12'd1219: coeff = 10'sd685;
		12'd1220: coeff = 10'sd686;
		12'd1221: coeff = 10'sd686;
		12'd1222: coeff = 10'sd687;
		12'd1223: coeff = 10'sd688;
		12'd1224: coeff = 10'sd689;
		12'd1225: coeff = 10'sd689;
		12'd1226: coeff = 10'sd690;
		12'd1227: coeff = 10'sd691;
		12'd1228: coeff = 10'sd692;
		12'd1229: coeff = 10'sd692;
		12'd1230: coeff = 10'sd693;
		12'd1231: coeff = 10'sd694;
		12'd1232: coeff = 10'sd695;
		12'd1233: coeff = 10'sd695;
		12'd1234: coeff = 10'sd696;
		12'd1235: coeff = 10'sd697;
		12'd1236: coeff = 10'sd698;
		12'd1237: coeff = 10'sd698;
		12'd1238: coeff = 10'sd699;
		12'd1239: coeff = 10'sd700;
		12'd1240: coeff = 10'sd701;
		12'd1241: coeff = 10'sd701;
		12'd1242: coeff = 10'sd702;
		12'd1243: coeff = 10'sd703;
		12'd1244: coeff = 10'sd704;
		12'd1245: coeff = 10'sd704;
		12'd1246: coeff = 10'sd705;
		12'd1247: coeff = 10'sd706;
		12'd1248: coeff = 10'sd707;
		12'd1249: coeff = 10'sd707;
		12'd1250: coeff = 10'sd708;
		12'd1251: coeff = 10'sd709;
		12'd1252: coeff = 10'sd710;
		12'd1253: coeff = 10'sd710;
		12'd1254: coeff = 10'sd711;
		12'd1255: coeff = 10'sd712;
		12'd1256: coeff = 10'sd713;
		12'd1257: coeff = 10'sd713;
		12'd1258: coeff = 10'sd714;
		12'd1259: coeff = 10'sd715;
		12'd1260: coeff = 10'sd716;
		12'd1261: coeff = 10'sd716;
		12'd1262: coeff = 10'sd717;
		12'd1263: coeff = 10'sd718;
		12'd1264: coeff = 10'sd719;
		12'd1265: coeff = 10'sd719;
		12'd1266: coeff = 10'sd720;
		12'd1267: coeff = 10'sd721;
		12'd1268: coeff = 10'sd721;
		12'd1269: coeff = 10'sd722;
		12'd1270: coeff = 10'sd723;
		12'd1271: coeff = 10'sd724;
		12'd1272: coeff = 10'sd724;
		12'd1273: coeff = 10'sd725;
		12'd1274: coeff = 10'sd726;
		12'd1275: coeff = 10'sd727;
		12'd1276: coeff = 10'sd727;
		12'd1277: coeff = 10'sd728;
		12'd1278: coeff = 10'sd729;
		12'd1279: coeff = 10'sd730;
		12'd1280: coeff = 10'sd730;
		12'd1281: coeff = 10'sd731;
		12'd1282: coeff = 10'sd732;
		12'd1283: coeff = 10'sd732;
		12'd1284: coeff = 10'sd733;
		12'd1285: coeff = 10'sd734;
		12'd1286: coeff = 10'sd735;
		12'd1287: coeff = 10'sd735;
		12'd1288: coeff = 10'sd736;
		12'd1289: coeff = 10'sd737;
		12'd1290: coeff = 10'sd737;
		12'd1291: coeff = 10'sd738;
		12'd1292: coeff = 10'sd739;
		12'd1293: coeff = 10'sd740;
		12'd1294: coeff = 10'sd740;
		12'd1295: coeff = 10'sd741;
		12'd1296: coeff = 10'sd742;
		12'd1297: coeff = 10'sd743;
		12'd1298: coeff = 10'sd743;
		12'd1299: coeff = 10'sd744;
		12'd1300: coeff = 10'sd745;
		12'd1301: coeff = 10'sd745;
		12'd1302: coeff = 10'sd746;
		12'd1303: coeff = 10'sd747;
		12'd1304: coeff = 10'sd748;
		12'd1305: coeff = 10'sd748;
		12'd1306: coeff = 10'sd749;
		12'd1307: coeff = 10'sd750;
		12'd1308: coeff = 10'sd750;
		12'd1309: coeff = 10'sd751;
		12'd1310: coeff = 10'sd752;
		12'd1311: coeff = 10'sd753;
		12'd1312: coeff = 10'sd753;
		12'd1313: coeff = 10'sd754;
		12'd1314: coeff = 10'sd755;
		12'd1315: coeff = 10'sd755;
		12'd1316: coeff = 10'sd756;
		12'd1317: coeff = 10'sd757;
		12'd1318: coeff = 10'sd757;
		12'd1319: coeff = 10'sd758;
		12'd1320: coeff = 10'sd759;
		12'd1321: coeff = 10'sd760;
		12'd1322: coeff = 10'sd760;
		12'd1323: coeff = 10'sd761;
		12'd1324: coeff = 10'sd762;
		12'd1325: coeff = 10'sd762;
		12'd1326: coeff = 10'sd763;
		12'd1327: coeff = 10'sd764;
		12'd1328: coeff = 10'sd765;
		12'd1329: coeff = 10'sd765;
		12'd1330: coeff = 10'sd766;
		12'd1331: coeff = 10'sd767;
		12'd1332: coeff = 10'sd767;
		12'd1333: coeff = 10'sd768;
		12'd1334: coeff = 10'sd769;
		12'd1335: coeff = 10'sd769;
		12'd1336: coeff = 10'sd770;
		12'd1337: coeff = 10'sd771;
		12'd1338: coeff = 10'sd771;
		12'd1339: coeff = 10'sd772;
		12'd1340: coeff = 10'sd773;
		12'd1341: coeff = 10'sd774;
		12'd1342: coeff = 10'sd774;
		12'd1343: coeff = 10'sd775;
		12'd1344: coeff = 10'sd776;
		12'd1345: coeff = 10'sd776;
		12'd1346: coeff = 10'sd777;
		12'd1347: coeff = 10'sd778;
		12'd1348: coeff = 10'sd778;
		12'd1349: coeff = 10'sd779;
		12'd1350: coeff = 10'sd780;
		12'd1351: coeff = 10'sd780;
		12'd1352: coeff = 10'sd781;
		12'd1353: coeff = 10'sd782;
		12'd1354: coeff = 10'sd782;
		12'd1355: coeff = 10'sd783;
		12'd1356: coeff = 10'sd784;
		12'd1357: coeff = 10'sd785;
		12'd1358: coeff = 10'sd785;
		12'd1359: coeff = 10'sd786;
		12'd1360: coeff = 10'sd787;
		12'd1361: coeff = 10'sd787;
		12'd1362: coeff = 10'sd788;
		12'd1363: coeff = 10'sd789;
		12'd1364: coeff = 10'sd789;
		12'd1365: coeff = 10'sd790;
		12'd1366: coeff = 10'sd791;
		12'd1367: coeff = 10'sd791;
		12'd1368: coeff = 10'sd792;
		12'd1369: coeff = 10'sd793;
		12'd1370: coeff = 10'sd793;
		12'd1371: coeff = 10'sd794;
		12'd1372: coeff = 10'sd795;
		12'd1373: coeff = 10'sd795;
		12'd1374: coeff = 10'sd796;
		12'd1375: coeff = 10'sd797;
		12'd1376: coeff = 10'sd797;
		12'd1377: coeff = 10'sd798;
		12'd1378: coeff = 10'sd799;
		12'd1379: coeff = 10'sd799;
		12'd1380: coeff = 10'sd800;
		12'd1381: coeff = 10'sd801;
		12'd1382: coeff = 10'sd801;
		12'd1383: coeff = 10'sd802;
		12'd1384: coeff = 10'sd803;
		12'd1385: coeff = 10'sd803;
		12'd1386: coeff = 10'sd804;
		12'd1387: coeff = 10'sd805;
		12'd1388: coeff = 10'sd805;
		12'd1389: coeff = 10'sd806;
		12'd1390: coeff = 10'sd807;
		12'd1391: coeff = 10'sd807;
		12'd1392: coeff = 10'sd808;
		12'd1393: coeff = 10'sd809;
		12'd1394: coeff = 10'sd809;
		12'd1395: coeff = 10'sd810;
		12'd1396: coeff = 10'sd811;
		12'd1397: coeff = 10'sd811;
		12'd1398: coeff = 10'sd812;
		12'd1399: coeff = 10'sd813;
		12'd1400: coeff = 10'sd813;
		12'd1401: coeff = 10'sd814;
		12'd1402: coeff = 10'sd814;
		12'd1403: coeff = 10'sd815;
		12'd1404: coeff = 10'sd816;
		12'd1405: coeff = 10'sd816;
		12'd1406: coeff = 10'sd817;
		12'd1407: coeff = 10'sd818;
		12'd1408: coeff = 10'sd818;
		12'd1409: coeff = 10'sd819;
		12'd1410: coeff = 10'sd820;
		12'd1411: coeff = 10'sd820;
		12'd1412: coeff = 10'sd821;
		12'd1413: coeff = 10'sd822;
		12'd1414: coeff = 10'sd822;
		12'd1415: coeff = 10'sd823;
		12'd1416: coeff = 10'sd823;
		12'd1417: coeff = 10'sd824;
		12'd1418: coeff = 10'sd825;
		12'd1419: coeff = 10'sd825;
		12'd1420: coeff = 10'sd826;
		12'd1421: coeff = 10'sd827;
		12'd1422: coeff = 10'sd827;
		12'd1423: coeff = 10'sd828;
		12'd1424: coeff = 10'sd829;
		12'd1425: coeff = 10'sd829;
		12'd1426: coeff = 10'sd830;
		12'd1427: coeff = 10'sd830;
		12'd1428: coeff = 10'sd831;
		12'd1429: coeff = 10'sd832;
		12'd1430: coeff = 10'sd832;
		12'd1431: coeff = 10'sd833;
		12'd1432: coeff = 10'sd834;
		12'd1433: coeff = 10'sd834;
		12'd1434: coeff = 10'sd835;
		12'd1435: coeff = 10'sd835;
		12'd1436: coeff = 10'sd836;
		12'd1437: coeff = 10'sd837;
		12'd1438: coeff = 10'sd837;
		12'd1439: coeff = 10'sd838;
		12'd1440: coeff = 10'sd839;
		12'd1441: coeff = 10'sd839;
		12'd1442: coeff = 10'sd840;
		12'd1443: coeff = 10'sd840;
		12'd1444: coeff = 10'sd841;
		12'd1445: coeff = 10'sd842;
		12'd1446: coeff = 10'sd842;
		12'd1447: coeff = 10'sd843;
		12'd1448: coeff = 10'sd844;
		12'd1449: coeff = 10'sd844;
		12'd1450: coeff = 10'sd845;
		12'd1451: coeff = 10'sd845;
		12'd1452: coeff = 10'sd846;
		12'd1453: coeff = 10'sd847;
		12'd1454: coeff = 10'sd847;
		12'd1455: coeff = 10'sd848;
		12'd1456: coeff = 10'sd848;
		12'd1457: coeff = 10'sd849;
		12'd1458: coeff = 10'sd850;
		12'd1459: coeff = 10'sd850;
		12'd1460: coeff = 10'sd851;
		12'd1461: coeff = 10'sd851;
		12'd1462: coeff = 10'sd852;
		12'd1463: coeff = 10'sd853;
		12'd1464: coeff = 10'sd853;
		12'd1465: coeff = 10'sd854;
		12'd1466: coeff = 10'sd854;
		12'd1467: coeff = 10'sd855;
		12'd1468: coeff = 10'sd856;
		12'd1469: coeff = 10'sd856;
		12'd1470: coeff = 10'sd857;
		12'd1471: coeff = 10'sd857;
		12'd1472: coeff = 10'sd858;
		12'd1473: coeff = 10'sd859;
		12'd1474: coeff = 10'sd859;
		12'd1475: coeff = 10'sd860;
		12'd1476: coeff = 10'sd860;
		12'd1477: coeff = 10'sd861;
		12'd1478: coeff = 10'sd862;
		12'd1479: coeff = 10'sd862;
		12'd1480: coeff = 10'sd863;
		12'd1481: coeff = 10'sd863;
		12'd1482: coeff = 10'sd864;
		12'd1483: coeff = 10'sd864;
		12'd1484: coeff = 10'sd865;
		12'd1485: coeff = 10'sd866;
		12'd1486: coeff = 10'sd866;
		12'd1487: coeff = 10'sd867;
		12'd1488: coeff = 10'sd867;
		12'd1489: coeff = 10'sd868;
		12'd1490: coeff = 10'sd869;
		12'd1491: coeff = 10'sd869;
		12'd1492: coeff = 10'sd870;
		12'd1493: coeff = 10'sd870;
		12'd1494: coeff = 10'sd871;
		12'd1495: coeff = 10'sd871;
		12'd1496: coeff = 10'sd872;
		12'd1497: coeff = 10'sd873;
		12'd1498: coeff = 10'sd873;
		12'd1499: coeff = 10'sd874;
		12'd1500: coeff = 10'sd874;
		12'd1501: coeff = 10'sd875;
		12'd1502: coeff = 10'sd875;
		12'd1503: coeff = 10'sd876;
		12'd1504: coeff = 10'sd877;
		12'd1505: coeff = 10'sd877;
		12'd1506: coeff = 10'sd878;
		12'd1507: coeff = 10'sd878;
		12'd1508: coeff = 10'sd879;
		12'd1509: coeff = 10'sd879;
		12'd1510: coeff = 10'sd880;
		12'd1511: coeff = 10'sd880;
		12'd1512: coeff = 10'sd881;
		12'd1513: coeff = 10'sd882;
		12'd1514: coeff = 10'sd882;
		12'd1515: coeff = 10'sd883;
		12'd1516: coeff = 10'sd883;
		12'd1517: coeff = 10'sd884;
		12'd1518: coeff = 10'sd884;
		12'd1519: coeff = 10'sd885;
		12'd1520: coeff = 10'sd885;
		12'd1521: coeff = 10'sd886;
		12'd1522: coeff = 10'sd887;
		12'd1523: coeff = 10'sd887;
		12'd1524: coeff = 10'sd888;
		12'd1525: coeff = 10'sd888;
		12'd1526: coeff = 10'sd889;
		12'd1527: coeff = 10'sd889;
		12'd1528: coeff = 10'sd890;
		12'd1529: coeff = 10'sd890;
		12'd1530: coeff = 10'sd891;
		12'd1531: coeff = 10'sd891;
		12'd1532: coeff = 10'sd892;
		12'd1533: coeff = 10'sd893;
		12'd1534: coeff = 10'sd893;
		12'd1535: coeff = 10'sd894;
		12'd1536: coeff = 10'sd894;
		12'd1537: coeff = 10'sd895;
		12'd1538: coeff = 10'sd895;
		12'd1539: coeff = 10'sd896;
		12'd1540: coeff = 10'sd896;
		12'd1541: coeff = 10'sd897;
		12'd1542: coeff = 10'sd897;
		12'd1543: coeff = 10'sd898;
		12'd1544: coeff = 10'sd898;
		12'd1545: coeff = 10'sd899;
		12'd1546: coeff = 10'sd899;
		12'd1547: coeff = 10'sd900;
		12'd1548: coeff = 10'sd900;
		12'd1549: coeff = 10'sd901;
		12'd1550: coeff = 10'sd902;
		12'd1551: coeff = 10'sd902;
		12'd1552: coeff = 10'sd903;
		12'd1553: coeff = 10'sd903;
		12'd1554: coeff = 10'sd904;
		12'd1555: coeff = 10'sd904;
		12'd1556: coeff = 10'sd905;
		12'd1557: coeff = 10'sd905;
		12'd1558: coeff = 10'sd906;
		12'd1559: coeff = 10'sd906;
		12'd1560: coeff = 10'sd907;
		12'd1561: coeff = 10'sd907;
		12'd1562: coeff = 10'sd908;
		12'd1563: coeff = 10'sd908;
		12'd1564: coeff = 10'sd909;
		12'd1565: coeff = 10'sd909;
		12'd1566: coeff = 10'sd910;
		12'd1567: coeff = 10'sd910;
		12'd1568: coeff = 10'sd911;
		12'd1569: coeff = 10'sd911;
		12'd1570: coeff = 10'sd912;
		12'd1571: coeff = 10'sd912;
		12'd1572: coeff = 10'sd913;
		12'd1573: coeff = 10'sd913;
		12'd1574: coeff = 10'sd914;
		12'd1575: coeff = 10'sd914;
		12'd1576: coeff = 10'sd915;
		12'd1577: coeff = 10'sd915;
		12'd1578: coeff = 10'sd916;
		12'd1579: coeff = 10'sd916;
		12'd1580: coeff = 10'sd917;
		12'd1581: coeff = 10'sd917;
		12'd1582: coeff = 10'sd918;
		12'd1583: coeff = 10'sd918;
		12'd1584: coeff = 10'sd919;
		12'd1585: coeff = 10'sd919;
		12'd1586: coeff = 10'sd920;
		12'd1587: coeff = 10'sd920;
		12'd1588: coeff = 10'sd921;
		12'd1589: coeff = 10'sd921;
		12'd1590: coeff = 10'sd922;
		12'd1591: coeff = 10'sd922;
		12'd1592: coeff = 10'sd923;
		12'd1593: coeff = 10'sd923;
		12'd1594: coeff = 10'sd924;
		12'd1595: coeff = 10'sd924;
		12'd1596: coeff = 10'sd925;
		12'd1597: coeff = 10'sd925;
		12'd1598: coeff = 10'sd925;
		12'd1599: coeff = 10'sd926;
		12'd1600: coeff = 10'sd926;
		12'd1601: coeff = 10'sd927;
		12'd1602: coeff = 10'sd927;
		12'd1603: coeff = 10'sd928;
		12'd1604: coeff = 10'sd928;
		12'd1605: coeff = 10'sd929;
		12'd1606: coeff = 10'sd929;
		12'd1607: coeff = 10'sd930;
		12'd1608: coeff = 10'sd930;
		12'd1609: coeff = 10'sd931;
		12'd1610: coeff = 10'sd931;
		12'd1611: coeff = 10'sd932;
		12'd1612: coeff = 10'sd932;
		12'd1613: coeff = 10'sd932;
		12'd1614: coeff = 10'sd933;
		12'd1615: coeff = 10'sd933;
		12'd1616: coeff = 10'sd934;
		12'd1617: coeff = 10'sd934;
		12'd1618: coeff = 10'sd935;
		12'd1619: coeff = 10'sd935;
		12'd1620: coeff = 10'sd936;
		12'd1621: coeff = 10'sd936;
		12'd1622: coeff = 10'sd937;
		12'd1623: coeff = 10'sd937;
		12'd1624: coeff = 10'sd937;
		12'd1625: coeff = 10'sd938;
		12'd1626: coeff = 10'sd938;
		12'd1627: coeff = 10'sd939;
		12'd1628: coeff = 10'sd939;
		12'd1629: coeff = 10'sd940;
		12'd1630: coeff = 10'sd940;
		12'd1631: coeff = 10'sd941;
		12'd1632: coeff = 10'sd941;
		12'd1633: coeff = 10'sd941;
		12'd1634: coeff = 10'sd942;
		12'd1635: coeff = 10'sd942;
		12'd1636: coeff = 10'sd943;
		12'd1637: coeff = 10'sd943;
		12'd1638: coeff = 10'sd944;
		12'd1639: coeff = 10'sd944;
		12'd1640: coeff = 10'sd944;
		12'd1641: coeff = 10'sd945;
		12'd1642: coeff = 10'sd945;
		12'd1643: coeff = 10'sd946;
		12'd1644: coeff = 10'sd946;
		12'd1645: coeff = 10'sd947;
		12'd1646: coeff = 10'sd947;
		12'd1647: coeff = 10'sd947;
		12'd1648: coeff = 10'sd948;
		12'd1649: coeff = 10'sd948;
		12'd1650: coeff = 10'sd949;
		12'd1651: coeff = 10'sd949;
		12'd1652: coeff = 10'sd950;
		12'd1653: coeff = 10'sd950;
		12'd1654: coeff = 10'sd950;
		12'd1655: coeff = 10'sd951;
		12'd1656: coeff = 10'sd951;
		12'd1657: coeff = 10'sd952;
		12'd1658: coeff = 10'sd952;
		12'd1659: coeff = 10'sd952;
		12'd1660: coeff = 10'sd953;
		12'd1661: coeff = 10'sd953;
		12'd1662: coeff = 10'sd954;
		12'd1663: coeff = 10'sd954;
		12'd1664: coeff = 10'sd954;
		12'd1665: coeff = 10'sd955;
		12'd1666: coeff = 10'sd955;
		12'd1667: coeff = 10'sd956;
		12'd1668: coeff = 10'sd956;
		12'd1669: coeff = 10'sd957;
		12'd1670: coeff = 10'sd957;
		12'd1671: coeff = 10'sd957;
		12'd1672: coeff = 10'sd958;
		12'd1673: coeff = 10'sd958;
		12'd1674: coeff = 10'sd958;
		12'd1675: coeff = 10'sd959;
		12'd1676: coeff = 10'sd959;
		12'd1677: coeff = 10'sd960;
		12'd1678: coeff = 10'sd960;
		12'd1679: coeff = 10'sd960;
		12'd1680: coeff = 10'sd961;
		12'd1681: coeff = 10'sd961;
		12'd1682: coeff = 10'sd962;
		12'd1683: coeff = 10'sd962;
		12'd1684: coeff = 10'sd962;
		12'd1685: coeff = 10'sd963;
		12'd1686: coeff = 10'sd963;
		12'd1687: coeff = 10'sd964;
		12'd1688: coeff = 10'sd964;
		12'd1689: coeff = 10'sd964;
		12'd1690: coeff = 10'sd965;
		12'd1691: coeff = 10'sd965;
		12'd1692: coeff = 10'sd965;
		12'd1693: coeff = 10'sd966;
		12'd1694: coeff = 10'sd966;
		12'd1695: coeff = 10'sd967;
		12'd1696: coeff = 10'sd967;
		12'd1697: coeff = 10'sd967;
		12'd1698: coeff = 10'sd968;
		12'd1699: coeff = 10'sd968;
		12'd1700: coeff = 10'sd968;
		12'd1701: coeff = 10'sd969;
		12'd1702: coeff = 10'sd969;
		12'd1703: coeff = 10'sd969;
		12'd1704: coeff = 10'sd970;
		12'd1705: coeff = 10'sd970;
		12'd1706: coeff = 10'sd971;
		12'd1707: coeff = 10'sd971;
		12'd1708: coeff = 10'sd971;
		12'd1709: coeff = 10'sd972;
		12'd1710: coeff = 10'sd972;
		12'd1711: coeff = 10'sd972;
		12'd1712: coeff = 10'sd973;
		12'd1713: coeff = 10'sd973;
		12'd1714: coeff = 10'sd973;
		12'd1715: coeff = 10'sd974;
		12'd1716: coeff = 10'sd974;
		12'd1717: coeff = 10'sd974;
		12'd1718: coeff = 10'sd975;
		12'd1719: coeff = 10'sd975;
		12'd1720: coeff = 10'sd975;
		12'd1721: coeff = 10'sd976;
		12'd1722: coeff = 10'sd976;
		12'd1723: coeff = 10'sd976;
		12'd1724: coeff = 10'sd977;
		12'd1725: coeff = 10'sd977;
		12'd1726: coeff = 10'sd977;
		12'd1727: coeff = 10'sd978;
		12'd1728: coeff = 10'sd978;
		12'd1729: coeff = 10'sd978;
		12'd1730: coeff = 10'sd979;
		12'd1731: coeff = 10'sd979;
		12'd1732: coeff = 10'sd979;
		12'd1733: coeff = 10'sd980;
		12'd1734: coeff = 10'sd980;
		12'd1735: coeff = 10'sd980;
		12'd1736: coeff = 10'sd981;
		12'd1737: coeff = 10'sd981;
		12'd1738: coeff = 10'sd981;
		12'd1739: coeff = 10'sd982;
		12'd1740: coeff = 10'sd982;
		12'd1741: coeff = 10'sd982;
		12'd1742: coeff = 10'sd983;
		12'd1743: coeff = 10'sd983;
		12'd1744: coeff = 10'sd983;
		12'd1745: coeff = 10'sd984;
		12'd1746: coeff = 10'sd984;
		12'd1747: coeff = 10'sd984;
		12'd1748: coeff = 10'sd985;
		12'd1749: coeff = 10'sd985;
		12'd1750: coeff = 10'sd985;
		12'd1751: coeff = 10'sd985;
		12'd1752: coeff = 10'sd986;
		12'd1753: coeff = 10'sd986;
		12'd1754: coeff = 10'sd986;
		12'd1755: coeff = 10'sd987;
		12'd1756: coeff = 10'sd987;
		12'd1757: coeff = 10'sd987;
		12'd1758: coeff = 10'sd988;
		12'd1759: coeff = 10'sd988;
		12'd1760: coeff = 10'sd988;
		12'd1761: coeff = 10'sd988;
		12'd1762: coeff = 10'sd989;
		12'd1763: coeff = 10'sd989;
		12'd1764: coeff = 10'sd989;
		12'd1765: coeff = 10'sd990;
		12'd1766: coeff = 10'sd990;
		12'd1767: coeff = 10'sd990;
		12'd1768: coeff = 10'sd991;
		12'd1769: coeff = 10'sd991;
		12'd1770: coeff = 10'sd991;
		12'd1771: coeff = 10'sd991;
		12'd1772: coeff = 10'sd992;
		12'd1773: coeff = 10'sd992;
		12'd1774: coeff = 10'sd992;
		12'd1775: coeff = 10'sd992;
		12'd1776: coeff = 10'sd993;
		12'd1777: coeff = 10'sd993;
		12'd1778: coeff = 10'sd993;
		12'd1779: coeff = 10'sd994;
		12'd1780: coeff = 10'sd994;
		12'd1781: coeff = 10'sd994;
		12'd1782: coeff = 10'sd994;
		12'd1783: coeff = 10'sd995;
		12'd1784: coeff = 10'sd995;
		12'd1785: coeff = 10'sd995;
		12'd1786: coeff = 10'sd995;
		12'd1787: coeff = 10'sd996;
		12'd1788: coeff = 10'sd996;
		12'd1789: coeff = 10'sd996;
		12'd1790: coeff = 10'sd997;
		12'd1791: coeff = 10'sd997;
		12'd1792: coeff = 10'sd997;
		12'd1793: coeff = 10'sd997;
		12'd1794: coeff = 10'sd998;
		12'd1795: coeff = 10'sd998;
		12'd1796: coeff = 10'sd998;
		12'd1797: coeff = 10'sd998;
		12'd1798: coeff = 10'sd999;
		12'd1799: coeff = 10'sd999;
		12'd1800: coeff = 10'sd999;
		12'd1801: coeff = 10'sd999;
		12'd1802: coeff = 10'sd1000;
		12'd1803: coeff = 10'sd1000;
		12'd1804: coeff = 10'sd1000;
		12'd1805: coeff = 10'sd1000;
		12'd1806: coeff = 10'sd1001;
		12'd1807: coeff = 10'sd1001;
		12'd1808: coeff = 10'sd1001;
		12'd1809: coeff = 10'sd1001;
		12'd1810: coeff = 10'sd1001;
		12'd1811: coeff = 10'sd1002;
		12'd1812: coeff = 10'sd1002;
		12'd1813: coeff = 10'sd1002;
		12'd1814: coeff = 10'sd1002;
		12'd1815: coeff = 10'sd1003;
		12'd1816: coeff = 10'sd1003;
		12'd1817: coeff = 10'sd1003;
		12'd1818: coeff = 10'sd1003;
		12'd1819: coeff = 10'sd1004;
		12'd1820: coeff = 10'sd1004;
		12'd1821: coeff = 10'sd1004;
		12'd1822: coeff = 10'sd1004;
		12'd1823: coeff = 10'sd1004;
		12'd1824: coeff = 10'sd1005;
		12'd1825: coeff = 10'sd1005;
		12'd1826: coeff = 10'sd1005;
		12'd1827: coeff = 10'sd1005;
		12'd1828: coeff = 10'sd1006;
		12'd1829: coeff = 10'sd1006;
		12'd1830: coeff = 10'sd1006;
		12'd1831: coeff = 10'sd1006;
		12'd1832: coeff = 10'sd1006;
		12'd1833: coeff = 10'sd1007;
		12'd1834: coeff = 10'sd1007;
		12'd1835: coeff = 10'sd1007;
		12'd1836: coeff = 10'sd1007;
		12'd1837: coeff = 10'sd1007;
		12'd1838: coeff = 10'sd1008;
		12'd1839: coeff = 10'sd1008;
		12'd1840: coeff = 10'sd1008;
		12'd1841: coeff = 10'sd1008;
		12'd1842: coeff = 10'sd1008;
		12'd1843: coeff = 10'sd1009;
		12'd1844: coeff = 10'sd1009;
		12'd1845: coeff = 10'sd1009;
		12'd1846: coeff = 10'sd1009;
		12'd1847: coeff = 10'sd1009;
		12'd1848: coeff = 10'sd1010;
		12'd1849: coeff = 10'sd1010;
		12'd1850: coeff = 10'sd1010;
		12'd1851: coeff = 10'sd1010;
		12'd1852: coeff = 10'sd1010;
		12'd1853: coeff = 10'sd1010;
		12'd1854: coeff = 10'sd1011;
		12'd1855: coeff = 10'sd1011;
		12'd1856: coeff = 10'sd1011;
		12'd1857: coeff = 10'sd1011;
		12'd1858: coeff = 10'sd1011;
		12'd1859: coeff = 10'sd1012;
		12'd1860: coeff = 10'sd1012;
		12'd1861: coeff = 10'sd1012;
		12'd1862: coeff = 10'sd1012;
		12'd1863: coeff = 10'sd1012;
		12'd1864: coeff = 10'sd1012;
		12'd1865: coeff = 10'sd1013;
		12'd1866: coeff = 10'sd1013;
		12'd1867: coeff = 10'sd1013;
		12'd1868: coeff = 10'sd1013;
		12'd1869: coeff = 10'sd1013;
		12'd1870: coeff = 10'sd1013;
		12'd1871: coeff = 10'sd1014;
		12'd1872: coeff = 10'sd1014;
		12'd1873: coeff = 10'sd1014;
		12'd1874: coeff = 10'sd1014;
		12'd1875: coeff = 10'sd1014;
		12'd1876: coeff = 10'sd1014;
		12'd1877: coeff = 10'sd1015;
		12'd1878: coeff = 10'sd1015;
		12'd1879: coeff = 10'sd1015;
		12'd1880: coeff = 10'sd1015;
		12'd1881: coeff = 10'sd1015;
		12'd1882: coeff = 10'sd1015;
		12'd1883: coeff = 10'sd1015;
		12'd1884: coeff = 10'sd1016;
		12'd1885: coeff = 10'sd1016;
		12'd1886: coeff = 10'sd1016;
		12'd1887: coeff = 10'sd1016;
		12'd1888: coeff = 10'sd1016;
		12'd1889: coeff = 10'sd1016;
		12'd1890: coeff = 10'sd1016;
		12'd1891: coeff = 10'sd1017;
		12'd1892: coeff = 10'sd1017;
		12'd1893: coeff = 10'sd1017;
		12'd1894: coeff = 10'sd1017;
		12'd1895: coeff = 10'sd1017;
		12'd1896: coeff = 10'sd1017;
		12'd1897: coeff = 10'sd1017;
		12'd1898: coeff = 10'sd1018;
		12'd1899: coeff = 10'sd1018;
		12'd1900: coeff = 10'sd1018;
		12'd1901: coeff = 10'sd1018;
		12'd1902: coeff = 10'sd1018;
		12'd1903: coeff = 10'sd1018;
		12'd1904: coeff = 10'sd1018;
		12'd1905: coeff = 10'sd1018;
		12'd1906: coeff = 10'sd1018;
		12'd1907: coeff = 10'sd1019;
		12'd1908: coeff = 10'sd1019;
		12'd1909: coeff = 10'sd1019;
		12'd1910: coeff = 10'sd1019;
		12'd1911: coeff = 10'sd1019;
		12'd1912: coeff = 10'sd1019;
		12'd1913: coeff = 10'sd1019;
		12'd1914: coeff = 10'sd1019;
		12'd1915: coeff = 10'sd1019;
		12'd1916: coeff = 10'sd1020;
		12'd1917: coeff = 10'sd1020;
		12'd1918: coeff = 10'sd1020;
		12'd1919: coeff = 10'sd1020;
		12'd1920: coeff = 10'sd1020;
		12'd1921: coeff = 10'sd1020;
		12'd1922: coeff = 10'sd1020;
		12'd1923: coeff = 10'sd1020;
		12'd1924: coeff = 10'sd1020;
		12'd1925: coeff = 10'sd1020;
		12'd1926: coeff = 10'sd1021;
		12'd1927: coeff = 10'sd1021;
		12'd1928: coeff = 10'sd1021;
		12'd1929: coeff = 10'sd1021;
		12'd1930: coeff = 10'sd1021;
		12'd1931: coeff = 10'sd1021;
		12'd1932: coeff = 10'sd1021;
		12'd1933: coeff = 10'sd1021;
		12'd1934: coeff = 10'sd1021;
		12'd1935: coeff = 10'sd1021;
		12'd1936: coeff = 10'sd1021;
		12'd1937: coeff = 10'sd1022;
		12'd1938: coeff = 10'sd1022;
		12'd1939: coeff = 10'sd1022;
		12'd1940: coeff = 10'sd1022;
		12'd1941: coeff = 10'sd1022;
		12'd1942: coeff = 10'sd1022;
		12'd1943: coeff = 10'sd1022;
		12'd1944: coeff = 10'sd1022;
		12'd1945: coeff = 10'sd1022;
		12'd1946: coeff = 10'sd1022;
		12'd1947: coeff = 10'sd1022;
		12'd1948: coeff = 10'sd1022;
		12'd1949: coeff = 10'sd1022;
		12'd1950: coeff = 10'sd1022;
		12'd1951: coeff = 10'sd1023;
		12'd1952: coeff = 10'sd1023;
		12'd1953: coeff = 10'sd1023;
		12'd1954: coeff = 10'sd1023;
		12'd1955: coeff = 10'sd1023;
		12'd1956: coeff = 10'sd1023;
		12'd1957: coeff = 10'sd1023;
		12'd1958: coeff = 10'sd1023;
		12'd1959: coeff = 10'sd1023;
		12'd1960: coeff = 10'sd1023;
		12'd1961: coeff = 10'sd1023;
		12'd1962: coeff = 10'sd1023;
		12'd1963: coeff = 10'sd1023;
		12'd1964: coeff = 10'sd1023;
		12'd1965: coeff = 10'sd1023;
		12'd1966: coeff = 10'sd1023;
		12'd1967: coeff = 10'sd1023;
		12'd1968: coeff = 10'sd1023;
		12'd1969: coeff = 10'sd1023;
		12'd1970: coeff = 10'sd1023;
		12'd1971: coeff = 10'sd1023;
		12'd1972: coeff = 10'sd1024;
		12'd1973: coeff = 10'sd1024;
		12'd1974: coeff = 10'sd1024;
		12'd1975: coeff = 10'sd1024;
		12'd1976: coeff = 10'sd1024;
		12'd1977: coeff = 10'sd1024;
		12'd1978: coeff = 10'sd1024;
		12'd1979: coeff = 10'sd1024;
		12'd1980: coeff = 10'sd1024;
		12'd1981: coeff = 10'sd1024;
		12'd1982: coeff = 10'sd1024;
		12'd1983: coeff = 10'sd1024;
		12'd1984: coeff = 10'sd1024;
		12'd1985: coeff = 10'sd1024;
		12'd1986: coeff = 10'sd1024;
		12'd1987: coeff = 10'sd1024;
		12'd1988: coeff = 10'sd1024;
		12'd1989: coeff = 10'sd1024;
		12'd1990: coeff = 10'sd1024;
		12'd1991: coeff = 10'sd1024;
		12'd1992: coeff = 10'sd1024;
		12'd1993: coeff = 10'sd1024;
		12'd1994: coeff = 10'sd1024;
		12'd1995: coeff = 10'sd1024;
		12'd1996: coeff = 10'sd1024;
		12'd1997: coeff = 10'sd1024;
		12'd1998: coeff = 10'sd1024;
		12'd1999: coeff = 10'sd1024;
		12'd2000: coeff = 10'sd1024;
		12'd2001: coeff = 10'sd1024;
		12'd2002: coeff = 10'sd1024;
		12'd2003: coeff = 10'sd1024;
		12'd2004: coeff = 10'sd1024;
		12'd2005: coeff = 10'sd1024;
		12'd2006: coeff = 10'sd1024;
		12'd2007: coeff = 10'sd1024;
		12'd2008: coeff = 10'sd1024;
		12'd2009: coeff = 10'sd1024;
		12'd2010: coeff = 10'sd1024;
		12'd2011: coeff = 10'sd1024;
		12'd2012: coeff = 10'sd1024;
		12'd2013: coeff = 10'sd1024;
		12'd2014: coeff = 10'sd1024;
		12'd2015: coeff = 10'sd1024;
		12'd2016: coeff = 10'sd1024;
		12'd2017: coeff = 10'sd1024;
		12'd2018: coeff = 10'sd1024;
		12'd2019: coeff = 10'sd1024;
		12'd2020: coeff = 10'sd1024;
		12'd2021: coeff = 10'sd1024;
		12'd2022: coeff = 10'sd1024;
		12'd2023: coeff = 10'sd1024;
		12'd2024: coeff = 10'sd1024;
		12'd2025: coeff = 10'sd1024;
		12'd2026: coeff = 10'sd1024;
		12'd2027: coeff = 10'sd1024;
		12'd2028: coeff = 10'sd1023;
		12'd2029: coeff = 10'sd1023;
		12'd2030: coeff = 10'sd1023;
		12'd2031: coeff = 10'sd1023;
		12'd2032: coeff = 10'sd1023;
		12'd2033: coeff = 10'sd1023;
		12'd2034: coeff = 10'sd1023;
		12'd2035: coeff = 10'sd1023;
		12'd2036: coeff = 10'sd1023;
		12'd2037: coeff = 10'sd1023;
		12'd2038: coeff = 10'sd1023;
		12'd2039: coeff = 10'sd1023;
		12'd2040: coeff = 10'sd1023;
		12'd2041: coeff = 10'sd1023;
		12'd2042: coeff = 10'sd1023;
		12'd2043: coeff = 10'sd1023;
		12'd2044: coeff = 10'sd1023;
		12'd2045: coeff = 10'sd1023;
		12'd2046: coeff = 10'sd1023;
		12'd2047: coeff = 10'sd1023;
		12'd2048: coeff = 10'sd1023;
		12'd2049: coeff = 10'sd1022;
		12'd2050: coeff = 10'sd1022;
		12'd2051: coeff = 10'sd1022;
		12'd2052: coeff = 10'sd1022;
		12'd2053: coeff = 10'sd1022;
		12'd2054: coeff = 10'sd1022;
		12'd2055: coeff = 10'sd1022;
		12'd2056: coeff = 10'sd1022;
		12'd2057: coeff = 10'sd1022;
		12'd2058: coeff = 10'sd1022;
		12'd2059: coeff = 10'sd1022;
		12'd2060: coeff = 10'sd1022;
		12'd2061: coeff = 10'sd1022;
		12'd2062: coeff = 10'sd1022;
		12'd2063: coeff = 10'sd1021;
		12'd2064: coeff = 10'sd1021;
		12'd2065: coeff = 10'sd1021;
		12'd2066: coeff = 10'sd1021;
		12'd2067: coeff = 10'sd1021;
		12'd2068: coeff = 10'sd1021;
		12'd2069: coeff = 10'sd1021;
		12'd2070: coeff = 10'sd1021;
		12'd2071: coeff = 10'sd1021;
		12'd2072: coeff = 10'sd1021;
		12'd2073: coeff = 10'sd1021;
		12'd2074: coeff = 10'sd1020;
		12'd2075: coeff = 10'sd1020;
		12'd2076: coeff = 10'sd1020;
		12'd2077: coeff = 10'sd1020;
		12'd2078: coeff = 10'sd1020;
		12'd2079: coeff = 10'sd1020;
		12'd2080: coeff = 10'sd1020;
		12'd2081: coeff = 10'sd1020;
		12'd2082: coeff = 10'sd1020;
		12'd2083: coeff = 10'sd1020;
		12'd2084: coeff = 10'sd1019;
		12'd2085: coeff = 10'sd1019;
		12'd2086: coeff = 10'sd1019;
		12'd2087: coeff = 10'sd1019;
		12'd2088: coeff = 10'sd1019;
		12'd2089: coeff = 10'sd1019;
		12'd2090: coeff = 10'sd1019;
		12'd2091: coeff = 10'sd1019;
		12'd2092: coeff = 10'sd1019;
		12'd2093: coeff = 10'sd1018;
		12'd2094: coeff = 10'sd1018;
		12'd2095: coeff = 10'sd1018;
		12'd2096: coeff = 10'sd1018;
		12'd2097: coeff = 10'sd1018;
		12'd2098: coeff = 10'sd1018;
		12'd2099: coeff = 10'sd1018;
		12'd2100: coeff = 10'sd1018;
		12'd2101: coeff = 10'sd1018;
		12'd2102: coeff = 10'sd1017;
		12'd2103: coeff = 10'sd1017;
		12'd2104: coeff = 10'sd1017;
		12'd2105: coeff = 10'sd1017;
		12'd2106: coeff = 10'sd1017;
		12'd2107: coeff = 10'sd1017;
		12'd2108: coeff = 10'sd1017;
		12'd2109: coeff = 10'sd1016;
		12'd2110: coeff = 10'sd1016;
		12'd2111: coeff = 10'sd1016;
		12'd2112: coeff = 10'sd1016;
		12'd2113: coeff = 10'sd1016;
		12'd2114: coeff = 10'sd1016;
		12'd2115: coeff = 10'sd1016;
		12'd2116: coeff = 10'sd1015;
		12'd2117: coeff = 10'sd1015;
		12'd2118: coeff = 10'sd1015;
		12'd2119: coeff = 10'sd1015;
		12'd2120: coeff = 10'sd1015;
		12'd2121: coeff = 10'sd1015;
		12'd2122: coeff = 10'sd1015;
		12'd2123: coeff = 10'sd1014;
		12'd2124: coeff = 10'sd1014;
		12'd2125: coeff = 10'sd1014;
		12'd2126: coeff = 10'sd1014;
		12'd2127: coeff = 10'sd1014;
		12'd2128: coeff = 10'sd1014;
		12'd2129: coeff = 10'sd1013;
		12'd2130: coeff = 10'sd1013;
		12'd2131: coeff = 10'sd1013;
		12'd2132: coeff = 10'sd1013;
		12'd2133: coeff = 10'sd1013;
		12'd2134: coeff = 10'sd1013;
		12'd2135: coeff = 10'sd1012;
		12'd2136: coeff = 10'sd1012;
		12'd2137: coeff = 10'sd1012;
		12'd2138: coeff = 10'sd1012;
		12'd2139: coeff = 10'sd1012;
		12'd2140: coeff = 10'sd1012;
		12'd2141: coeff = 10'sd1011;
		12'd2142: coeff = 10'sd1011;
		12'd2143: coeff = 10'sd1011;
		12'd2144: coeff = 10'sd1011;
		12'd2145: coeff = 10'sd1011;
		12'd2146: coeff = 10'sd1010;
		12'd2147: coeff = 10'sd1010;
		12'd2148: coeff = 10'sd1010;
		12'd2149: coeff = 10'sd1010;
		12'd2150: coeff = 10'sd1010;
		12'd2151: coeff = 10'sd1010;
		12'd2152: coeff = 10'sd1009;
		12'd2153: coeff = 10'sd1009;
		12'd2154: coeff = 10'sd1009;
		12'd2155: coeff = 10'sd1009;
		12'd2156: coeff = 10'sd1009;
		12'd2157: coeff = 10'sd1008;
		12'd2158: coeff = 10'sd1008;
		12'd2159: coeff = 10'sd1008;
		12'd2160: coeff = 10'sd1008;
		12'd2161: coeff = 10'sd1008;
		12'd2162: coeff = 10'sd1007;
		12'd2163: coeff = 10'sd1007;
		12'd2164: coeff = 10'sd1007;
		12'd2165: coeff = 10'sd1007;
		12'd2166: coeff = 10'sd1007;
		12'd2167: coeff = 10'sd1006;
		12'd2168: coeff = 10'sd1006;
		12'd2169: coeff = 10'sd1006;
		12'd2170: coeff = 10'sd1006;
		12'd2171: coeff = 10'sd1006;
		12'd2172: coeff = 10'sd1005;
		12'd2173: coeff = 10'sd1005;
		12'd2174: coeff = 10'sd1005;
		12'd2175: coeff = 10'sd1005;
		12'd2176: coeff = 10'sd1004;
		12'd2177: coeff = 10'sd1004;
		12'd2178: coeff = 10'sd1004;
		12'd2179: coeff = 10'sd1004;
		12'd2180: coeff = 10'sd1004;
		12'd2181: coeff = 10'sd1003;
		12'd2182: coeff = 10'sd1003;
		12'd2183: coeff = 10'sd1003;
		12'd2184: coeff = 10'sd1003;
		12'd2185: coeff = 10'sd1002;
		12'd2186: coeff = 10'sd1002;
		12'd2187: coeff = 10'sd1002;
		12'd2188: coeff = 10'sd1002;
		12'd2189: coeff = 10'sd1001;
		12'd2190: coeff = 10'sd1001;
		12'd2191: coeff = 10'sd1001;
		12'd2192: coeff = 10'sd1001;
		12'd2193: coeff = 10'sd1001;
		12'd2194: coeff = 10'sd1000;
		12'd2195: coeff = 10'sd1000;
		12'd2196: coeff = 10'sd1000;
		12'd2197: coeff = 10'sd1000;
		12'd2198: coeff = 10'sd999;
		12'd2199: coeff = 10'sd999;
		12'd2200: coeff = 10'sd999;
		12'd2201: coeff = 10'sd999;
		12'd2202: coeff = 10'sd998;
		12'd2203: coeff = 10'sd998;
		12'd2204: coeff = 10'sd998;
		12'd2205: coeff = 10'sd998;
		12'd2206: coeff = 10'sd997;
		12'd2207: coeff = 10'sd997;
		12'd2208: coeff = 10'sd997;
		12'd2209: coeff = 10'sd997;
		12'd2210: coeff = 10'sd996;
		12'd2211: coeff = 10'sd996;
		12'd2212: coeff = 10'sd996;
		12'd2213: coeff = 10'sd995;
		12'd2214: coeff = 10'sd995;
		12'd2215: coeff = 10'sd995;
		12'd2216: coeff = 10'sd995;
		12'd2217: coeff = 10'sd994;
		12'd2218: coeff = 10'sd994;
		12'd2219: coeff = 10'sd994;
		12'd2220: coeff = 10'sd994;
		12'd2221: coeff = 10'sd993;
		12'd2222: coeff = 10'sd993;
		12'd2223: coeff = 10'sd993;
		12'd2224: coeff = 10'sd992;
		12'd2225: coeff = 10'sd992;
		12'd2226: coeff = 10'sd992;
		12'd2227: coeff = 10'sd992;
		12'd2228: coeff = 10'sd991;
		12'd2229: coeff = 10'sd991;
		12'd2230: coeff = 10'sd991;
		12'd2231: coeff = 10'sd991;
		12'd2232: coeff = 10'sd990;
		12'd2233: coeff = 10'sd990;
		12'd2234: coeff = 10'sd990;
		12'd2235: coeff = 10'sd989;
		12'd2236: coeff = 10'sd989;
		12'd2237: coeff = 10'sd989;
		12'd2238: coeff = 10'sd988;
		12'd2239: coeff = 10'sd988;
		12'd2240: coeff = 10'sd988;
		12'd2241: coeff = 10'sd988;
		12'd2242: coeff = 10'sd987;
		12'd2243: coeff = 10'sd987;
		12'd2244: coeff = 10'sd987;
		12'd2245: coeff = 10'sd986;
		12'd2246: coeff = 10'sd986;
		12'd2247: coeff = 10'sd986;
		12'd2248: coeff = 10'sd985;
		12'd2249: coeff = 10'sd985;
		12'd2250: coeff = 10'sd985;
		12'd2251: coeff = 10'sd985;
		12'd2252: coeff = 10'sd984;
		12'd2253: coeff = 10'sd984;
		12'd2254: coeff = 10'sd984;
		12'd2255: coeff = 10'sd983;
		12'd2256: coeff = 10'sd983;
		12'd2257: coeff = 10'sd983;
		12'd2258: coeff = 10'sd982;
		12'd2259: coeff = 10'sd982;
		12'd2260: coeff = 10'sd982;
		12'd2261: coeff = 10'sd981;
		12'd2262: coeff = 10'sd981;
		12'd2263: coeff = 10'sd981;
		12'd2264: coeff = 10'sd980;
		12'd2265: coeff = 10'sd980;
		12'd2266: coeff = 10'sd980;
		12'd2267: coeff = 10'sd979;
		12'd2268: coeff = 10'sd979;
		12'd2269: coeff = 10'sd979;
		12'd2270: coeff = 10'sd978;
		12'd2271: coeff = 10'sd978;
		12'd2272: coeff = 10'sd978;
		12'd2273: coeff = 10'sd977;
		12'd2274: coeff = 10'sd977;
		12'd2275: coeff = 10'sd977;
		12'd2276: coeff = 10'sd976;
		12'd2277: coeff = 10'sd976;
		12'd2278: coeff = 10'sd976;
		12'd2279: coeff = 10'sd975;
		12'd2280: coeff = 10'sd975;
		12'd2281: coeff = 10'sd975;
		12'd2282: coeff = 10'sd974;
		12'd2283: coeff = 10'sd974;
		12'd2284: coeff = 10'sd974;
		12'd2285: coeff = 10'sd973;
		12'd2286: coeff = 10'sd973;
		12'd2287: coeff = 10'sd973;
		12'd2288: coeff = 10'sd972;
		12'd2289: coeff = 10'sd972;
		12'd2290: coeff = 10'sd972;
		12'd2291: coeff = 10'sd971;
		12'd2292: coeff = 10'sd971;
		12'd2293: coeff = 10'sd971;
		12'd2294: coeff = 10'sd970;
		12'd2295: coeff = 10'sd970;
		12'd2296: coeff = 10'sd969;
		12'd2297: coeff = 10'sd969;
		12'd2298: coeff = 10'sd969;
		12'd2299: coeff = 10'sd968;
		12'd2300: coeff = 10'sd968;
		12'd2301: coeff = 10'sd968;
		12'd2302: coeff = 10'sd967;
		12'd2303: coeff = 10'sd967;
		12'd2304: coeff = 10'sd967;
		12'd2305: coeff = 10'sd966;
		12'd2306: coeff = 10'sd966;
		12'd2307: coeff = 10'sd965;
		12'd2308: coeff = 10'sd965;
		12'd2309: coeff = 10'sd965;
		12'd2310: coeff = 10'sd964;
		12'd2311: coeff = 10'sd964;
		12'd2312: coeff = 10'sd964;
		12'd2313: coeff = 10'sd963;
		12'd2314: coeff = 10'sd963;
		12'd2315: coeff = 10'sd962;
		12'd2316: coeff = 10'sd962;
		12'd2317: coeff = 10'sd962;
		12'd2318: coeff = 10'sd961;
		12'd2319: coeff = 10'sd961;
		12'd2320: coeff = 10'sd960;
		12'd2321: coeff = 10'sd960;
		12'd2322: coeff = 10'sd960;
		12'd2323: coeff = 10'sd959;
		12'd2324: coeff = 10'sd959;
		12'd2325: coeff = 10'sd958;
		12'd2326: coeff = 10'sd958;
		12'd2327: coeff = 10'sd958;
		12'd2328: coeff = 10'sd957;
		12'd2329: coeff = 10'sd957;
		12'd2330: coeff = 10'sd957;
		12'd2331: coeff = 10'sd956;
		12'd2332: coeff = 10'sd956;
		12'd2333: coeff = 10'sd955;
		12'd2334: coeff = 10'sd955;
		12'd2335: coeff = 10'sd954;
		12'd2336: coeff = 10'sd954;
		12'd2337: coeff = 10'sd954;
		12'd2338: coeff = 10'sd953;
		12'd2339: coeff = 10'sd953;
		12'd2340: coeff = 10'sd952;
		12'd2341: coeff = 10'sd952;
		12'd2342: coeff = 10'sd952;
		12'd2343: coeff = 10'sd951;
		12'd2344: coeff = 10'sd951;
		12'd2345: coeff = 10'sd950;
		12'd2346: coeff = 10'sd950;
		12'd2347: coeff = 10'sd950;
		12'd2348: coeff = 10'sd949;
		12'd2349: coeff = 10'sd949;
		12'd2350: coeff = 10'sd948;
		12'd2351: coeff = 10'sd948;
		12'd2352: coeff = 10'sd947;
		12'd2353: coeff = 10'sd947;
		12'd2354: coeff = 10'sd947;
		12'd2355: coeff = 10'sd946;
		12'd2356: coeff = 10'sd946;
		12'd2357: coeff = 10'sd945;
		12'd2358: coeff = 10'sd945;
		12'd2359: coeff = 10'sd944;
		12'd2360: coeff = 10'sd944;
		12'd2361: coeff = 10'sd944;
		12'd2362: coeff = 10'sd943;
		12'd2363: coeff = 10'sd943;
		12'd2364: coeff = 10'sd942;
		12'd2365: coeff = 10'sd942;
		12'd2366: coeff = 10'sd941;
		12'd2367: coeff = 10'sd941;
		12'd2368: coeff = 10'sd941;
		12'd2369: coeff = 10'sd940;
		12'd2370: coeff = 10'sd940;
		12'd2371: coeff = 10'sd939;
		12'd2372: coeff = 10'sd939;
		12'd2373: coeff = 10'sd938;
		12'd2374: coeff = 10'sd938;
		12'd2375: coeff = 10'sd937;
		12'd2376: coeff = 10'sd937;
		12'd2377: coeff = 10'sd937;
		12'd2378: coeff = 10'sd936;
		12'd2379: coeff = 10'sd936;
		12'd2380: coeff = 10'sd935;
		12'd2381: coeff = 10'sd935;
		12'd2382: coeff = 10'sd934;
		12'd2383: coeff = 10'sd934;
		12'd2384: coeff = 10'sd933;
		12'd2385: coeff = 10'sd933;
		12'd2386: coeff = 10'sd932;
		12'd2387: coeff = 10'sd932;
		12'd2388: coeff = 10'sd932;
		12'd2389: coeff = 10'sd931;
		12'd2390: coeff = 10'sd931;
		12'd2391: coeff = 10'sd930;
		12'd2392: coeff = 10'sd930;
		12'd2393: coeff = 10'sd929;
		12'd2394: coeff = 10'sd929;
		12'd2395: coeff = 10'sd928;
		12'd2396: coeff = 10'sd928;
		12'd2397: coeff = 10'sd927;
		12'd2398: coeff = 10'sd927;
		12'd2399: coeff = 10'sd926;
		12'd2400: coeff = 10'sd926;
		12'd2401: coeff = 10'sd925;
		12'd2402: coeff = 10'sd925;
		12'd2403: coeff = 10'sd925;
		12'd2404: coeff = 10'sd924;
		12'd2405: coeff = 10'sd924;
		12'd2406: coeff = 10'sd923;
		12'd2407: coeff = 10'sd923;
		12'd2408: coeff = 10'sd922;
		12'd2409: coeff = 10'sd922;
		12'd2410: coeff = 10'sd921;
		12'd2411: coeff = 10'sd921;
		12'd2412: coeff = 10'sd920;
		12'd2413: coeff = 10'sd920;
		12'd2414: coeff = 10'sd919;
		12'd2415: coeff = 10'sd919;
		12'd2416: coeff = 10'sd918;
		12'd2417: coeff = 10'sd918;
		12'd2418: coeff = 10'sd917;
		12'd2419: coeff = 10'sd917;
		12'd2420: coeff = 10'sd916;
		12'd2421: coeff = 10'sd916;
		12'd2422: coeff = 10'sd915;
		12'd2423: coeff = 10'sd915;
		12'd2424: coeff = 10'sd914;
		12'd2425: coeff = 10'sd914;
		12'd2426: coeff = 10'sd913;
		12'd2427: coeff = 10'sd913;
		12'd2428: coeff = 10'sd912;
		12'd2429: coeff = 10'sd912;
		12'd2430: coeff = 10'sd911;
		12'd2431: coeff = 10'sd911;
		12'd2432: coeff = 10'sd910;
		12'd2433: coeff = 10'sd910;
		12'd2434: coeff = 10'sd909;
		12'd2435: coeff = 10'sd909;
		12'd2436: coeff = 10'sd908;
		12'd2437: coeff = 10'sd908;
		12'd2438: coeff = 10'sd907;
		12'd2439: coeff = 10'sd907;
		12'd2440: coeff = 10'sd906;
		12'd2441: coeff = 10'sd906;
		12'd2442: coeff = 10'sd905;
		12'd2443: coeff = 10'sd905;
		12'd2444: coeff = 10'sd904;
		12'd2445: coeff = 10'sd904;
		12'd2446: coeff = 10'sd903;
		12'd2447: coeff = 10'sd903;
		12'd2448: coeff = 10'sd902;
		12'd2449: coeff = 10'sd902;
		12'd2450: coeff = 10'sd901;
		12'd2451: coeff = 10'sd900;
		12'd2452: coeff = 10'sd900;
		12'd2453: coeff = 10'sd899;
		12'd2454: coeff = 10'sd899;
		12'd2455: coeff = 10'sd898;
		12'd2456: coeff = 10'sd898;
		12'd2457: coeff = 10'sd897;
		12'd2458: coeff = 10'sd897;
		12'd2459: coeff = 10'sd896;
		12'd2460: coeff = 10'sd896;
		12'd2461: coeff = 10'sd895;
		12'd2462: coeff = 10'sd895;
		12'd2463: coeff = 10'sd894;
		12'd2464: coeff = 10'sd894;
		12'd2465: coeff = 10'sd893;
		12'd2466: coeff = 10'sd893;
		12'd2467: coeff = 10'sd892;
		12'd2468: coeff = 10'sd891;
		12'd2469: coeff = 10'sd891;
		12'd2470: coeff = 10'sd890;
		12'd2471: coeff = 10'sd890;
		12'd2472: coeff = 10'sd889;
		12'd2473: coeff = 10'sd889;
		12'd2474: coeff = 10'sd888;
		12'd2475: coeff = 10'sd888;
		12'd2476: coeff = 10'sd887;
		12'd2477: coeff = 10'sd887;
		12'd2478: coeff = 10'sd886;
		12'd2479: coeff = 10'sd885;
		12'd2480: coeff = 10'sd885;
		12'd2481: coeff = 10'sd884;
		12'd2482: coeff = 10'sd884;
		12'd2483: coeff = 10'sd883;
		12'd2484: coeff = 10'sd883;
		12'd2485: coeff = 10'sd882;
		12'd2486: coeff = 10'sd882;
		12'd2487: coeff = 10'sd881;
		12'd2488: coeff = 10'sd880;
		12'd2489: coeff = 10'sd880;
		12'd2490: coeff = 10'sd879;
		12'd2491: coeff = 10'sd879;
		12'd2492: coeff = 10'sd878;
		12'd2493: coeff = 10'sd878;
		12'd2494: coeff = 10'sd877;
		12'd2495: coeff = 10'sd877;
		12'd2496: coeff = 10'sd876;
		12'd2497: coeff = 10'sd875;
		12'd2498: coeff = 10'sd875;
		12'd2499: coeff = 10'sd874;
		12'd2500: coeff = 10'sd874;
		12'd2501: coeff = 10'sd873;
		12'd2502: coeff = 10'sd873;
		12'd2503: coeff = 10'sd872;
		12'd2504: coeff = 10'sd871;
		12'd2505: coeff = 10'sd871;
		12'd2506: coeff = 10'sd870;
		12'd2507: coeff = 10'sd870;
		12'd2508: coeff = 10'sd869;
		12'd2509: coeff = 10'sd869;
		12'd2510: coeff = 10'sd868;
		12'd2511: coeff = 10'sd867;
		12'd2512: coeff = 10'sd867;
		12'd2513: coeff = 10'sd866;
		12'd2514: coeff = 10'sd866;
		12'd2515: coeff = 10'sd865;
		12'd2516: coeff = 10'sd864;
		12'd2517: coeff = 10'sd864;
		12'd2518: coeff = 10'sd863;
		12'd2519: coeff = 10'sd863;
		12'd2520: coeff = 10'sd862;
		12'd2521: coeff = 10'sd862;
		12'd2522: coeff = 10'sd861;
		12'd2523: coeff = 10'sd860;
		12'd2524: coeff = 10'sd860;
		12'd2525: coeff = 10'sd859;
		12'd2526: coeff = 10'sd859;
		12'd2527: coeff = 10'sd858;
		12'd2528: coeff = 10'sd857;
		12'd2529: coeff = 10'sd857;
		12'd2530: coeff = 10'sd856;
		12'd2531: coeff = 10'sd856;
		12'd2532: coeff = 10'sd855;
		12'd2533: coeff = 10'sd854;
		12'd2534: coeff = 10'sd854;
		12'd2535: coeff = 10'sd853;
		12'd2536: coeff = 10'sd853;
		12'd2537: coeff = 10'sd852;
		12'd2538: coeff = 10'sd851;
		12'd2539: coeff = 10'sd851;
		12'd2540: coeff = 10'sd850;
		12'd2541: coeff = 10'sd850;
		12'd2542: coeff = 10'sd849;
		12'd2543: coeff = 10'sd848;
		12'd2544: coeff = 10'sd848;
		12'd2545: coeff = 10'sd847;
		12'd2546: coeff = 10'sd847;
		12'd2547: coeff = 10'sd846;
		12'd2548: coeff = 10'sd845;
		12'd2549: coeff = 10'sd845;
		12'd2550: coeff = 10'sd844;
		12'd2551: coeff = 10'sd844;
		12'd2552: coeff = 10'sd843;
		12'd2553: coeff = 10'sd842;
		12'd2554: coeff = 10'sd842;
		12'd2555: coeff = 10'sd841;
		12'd2556: coeff = 10'sd840;
		12'd2557: coeff = 10'sd840;
		12'd2558: coeff = 10'sd839;
		12'd2559: coeff = 10'sd839;
		12'd2560: coeff = 10'sd838;
		12'd2561: coeff = 10'sd837;
		12'd2562: coeff = 10'sd837;
		12'd2563: coeff = 10'sd836;
		12'd2564: coeff = 10'sd835;
		12'd2565: coeff = 10'sd835;
		12'd2566: coeff = 10'sd834;
		12'd2567: coeff = 10'sd834;
		12'd2568: coeff = 10'sd833;
		12'd2569: coeff = 10'sd832;
		12'd2570: coeff = 10'sd832;
		12'd2571: coeff = 10'sd831;
		12'd2572: coeff = 10'sd830;
		12'd2573: coeff = 10'sd830;
		12'd2574: coeff = 10'sd829;
		12'd2575: coeff = 10'sd829;
		12'd2576: coeff = 10'sd828;
		12'd2577: coeff = 10'sd827;
		12'd2578: coeff = 10'sd827;
		12'd2579: coeff = 10'sd826;
		12'd2580: coeff = 10'sd825;
		12'd2581: coeff = 10'sd825;
		12'd2582: coeff = 10'sd824;
		12'd2583: coeff = 10'sd823;
		12'd2584: coeff = 10'sd823;
		12'd2585: coeff = 10'sd822;
		12'd2586: coeff = 10'sd822;
		12'd2587: coeff = 10'sd821;
		12'd2588: coeff = 10'sd820;
		12'd2589: coeff = 10'sd820;
		12'd2590: coeff = 10'sd819;
		12'd2591: coeff = 10'sd818;
		12'd2592: coeff = 10'sd818;
		12'd2593: coeff = 10'sd817;
		12'd2594: coeff = 10'sd816;
		12'd2595: coeff = 10'sd816;
		12'd2596: coeff = 10'sd815;
		12'd2597: coeff = 10'sd814;
		12'd2598: coeff = 10'sd814;
		12'd2599: coeff = 10'sd813;
		12'd2600: coeff = 10'sd813;
		12'd2601: coeff = 10'sd812;
		12'd2602: coeff = 10'sd811;
		12'd2603: coeff = 10'sd811;
		12'd2604: coeff = 10'sd810;
		12'd2605: coeff = 10'sd809;
		12'd2606: coeff = 10'sd809;
		12'd2607: coeff = 10'sd808;
		12'd2608: coeff = 10'sd807;
		12'd2609: coeff = 10'sd807;
		12'd2610: coeff = 10'sd806;
		12'd2611: coeff = 10'sd805;
		12'd2612: coeff = 10'sd805;
		12'd2613: coeff = 10'sd804;
		12'd2614: coeff = 10'sd803;
		12'd2615: coeff = 10'sd803;
		12'd2616: coeff = 10'sd802;
		12'd2617: coeff = 10'sd801;
		12'd2618: coeff = 10'sd801;
		12'd2619: coeff = 10'sd800;
		12'd2620: coeff = 10'sd799;
		12'd2621: coeff = 10'sd799;
		12'd2622: coeff = 10'sd798;
		12'd2623: coeff = 10'sd797;
		12'd2624: coeff = 10'sd797;
		12'd2625: coeff = 10'sd796;
		12'd2626: coeff = 10'sd795;
		12'd2627: coeff = 10'sd795;
		12'd2628: coeff = 10'sd794;
		12'd2629: coeff = 10'sd793;
		12'd2630: coeff = 10'sd793;
		12'd2631: coeff = 10'sd792;
		12'd2632: coeff = 10'sd791;
		12'd2633: coeff = 10'sd791;
		12'd2634: coeff = 10'sd790;
		12'd2635: coeff = 10'sd789;
		12'd2636: coeff = 10'sd789;
		12'd2637: coeff = 10'sd788;
		12'd2638: coeff = 10'sd787;
		12'd2639: coeff = 10'sd787;
		12'd2640: coeff = 10'sd786;
		12'd2641: coeff = 10'sd785;
		12'd2642: coeff = 10'sd785;
		12'd2643: coeff = 10'sd784;
		12'd2644: coeff = 10'sd783;
		12'd2645: coeff = 10'sd782;
		12'd2646: coeff = 10'sd782;
		12'd2647: coeff = 10'sd781;
		12'd2648: coeff = 10'sd780;
		12'd2649: coeff = 10'sd780;
		12'd2650: coeff = 10'sd779;
		12'd2651: coeff = 10'sd778;
		12'd2652: coeff = 10'sd778;
		12'd2653: coeff = 10'sd777;
		12'd2654: coeff = 10'sd776;
		12'd2655: coeff = 10'sd776;
		12'd2656: coeff = 10'sd775;
		12'd2657: coeff = 10'sd774;
		12'd2658: coeff = 10'sd774;
		12'd2659: coeff = 10'sd773;
		12'd2660: coeff = 10'sd772;
		12'd2661: coeff = 10'sd771;
		12'd2662: coeff = 10'sd771;
		12'd2663: coeff = 10'sd770;
		12'd2664: coeff = 10'sd769;
		12'd2665: coeff = 10'sd769;
		12'd2666: coeff = 10'sd768;
		12'd2667: coeff = 10'sd767;
		12'd2668: coeff = 10'sd767;
		12'd2669: coeff = 10'sd766;
		12'd2670: coeff = 10'sd765;
		12'd2671: coeff = 10'sd765;
		12'd2672: coeff = 10'sd764;
		12'd2673: coeff = 10'sd763;
		12'd2674: coeff = 10'sd762;
		12'd2675: coeff = 10'sd762;
		12'd2676: coeff = 10'sd761;
		12'd2677: coeff = 10'sd760;
		12'd2678: coeff = 10'sd760;
		12'd2679: coeff = 10'sd759;
		12'd2680: coeff = 10'sd758;
		12'd2681: coeff = 10'sd757;
		12'd2682: coeff = 10'sd757;
		12'd2683: coeff = 10'sd756;
		12'd2684: coeff = 10'sd755;
		12'd2685: coeff = 10'sd755;
		12'd2686: coeff = 10'sd754;
		12'd2687: coeff = 10'sd753;
		12'd2688: coeff = 10'sd753;
		12'd2689: coeff = 10'sd752;
		12'd2690: coeff = 10'sd751;
		12'd2691: coeff = 10'sd750;
		12'd2692: coeff = 10'sd750;
		12'd2693: coeff = 10'sd749;
		12'd2694: coeff = 10'sd748;
		12'd2695: coeff = 10'sd748;
		12'd2696: coeff = 10'sd747;
		12'd2697: coeff = 10'sd746;
		12'd2698: coeff = 10'sd745;
		12'd2699: coeff = 10'sd745;
		12'd2700: coeff = 10'sd744;
		12'd2701: coeff = 10'sd743;
		12'd2702: coeff = 10'sd743;
		12'd2703: coeff = 10'sd742;
		12'd2704: coeff = 10'sd741;
		12'd2705: coeff = 10'sd740;
		12'd2706: coeff = 10'sd740;
		12'd2707: coeff = 10'sd739;
		12'd2708: coeff = 10'sd738;
		12'd2709: coeff = 10'sd737;
		12'd2710: coeff = 10'sd737;
		12'd2711: coeff = 10'sd736;
		12'd2712: coeff = 10'sd735;
		12'd2713: coeff = 10'sd735;
		12'd2714: coeff = 10'sd734;
		12'd2715: coeff = 10'sd733;
		12'd2716: coeff = 10'sd732;
		12'd2717: coeff = 10'sd732;
		12'd2718: coeff = 10'sd731;
		12'd2719: coeff = 10'sd730;
		12'd2720: coeff = 10'sd730;
		12'd2721: coeff = 10'sd729;
		12'd2722: coeff = 10'sd728;
		12'd2723: coeff = 10'sd727;
		12'd2724: coeff = 10'sd727;
		12'd2725: coeff = 10'sd726;
		12'd2726: coeff = 10'sd725;
		12'd2727: coeff = 10'sd724;
		12'd2728: coeff = 10'sd724;
		12'd2729: coeff = 10'sd723;
		12'd2730: coeff = 10'sd722;
		12'd2731: coeff = 10'sd721;
		12'd2732: coeff = 10'sd721;
		12'd2733: coeff = 10'sd720;
		12'd2734: coeff = 10'sd719;
		12'd2735: coeff = 10'sd719;
		12'd2736: coeff = 10'sd718;
		12'd2737: coeff = 10'sd717;
		12'd2738: coeff = 10'sd716;
		12'd2739: coeff = 10'sd716;
		12'd2740: coeff = 10'sd715;
		12'd2741: coeff = 10'sd714;
		12'd2742: coeff = 10'sd713;
		12'd2743: coeff = 10'sd713;
		12'd2744: coeff = 10'sd712;
		12'd2745: coeff = 10'sd711;
		12'd2746: coeff = 10'sd710;
		12'd2747: coeff = 10'sd710;
		12'd2748: coeff = 10'sd709;
		12'd2749: coeff = 10'sd708;
		12'd2750: coeff = 10'sd707;
		12'd2751: coeff = 10'sd707;
		12'd2752: coeff = 10'sd706;
		12'd2753: coeff = 10'sd705;
		12'd2754: coeff = 10'sd704;
		12'd2755: coeff = 10'sd704;
		12'd2756: coeff = 10'sd703;
		12'd2757: coeff = 10'sd702;
		12'd2758: coeff = 10'sd701;
		12'd2759: coeff = 10'sd701;
		12'd2760: coeff = 10'sd700;
		12'd2761: coeff = 10'sd699;
		12'd2762: coeff = 10'sd698;
		12'd2763: coeff = 10'sd698;
		12'd2764: coeff = 10'sd697;
		12'd2765: coeff = 10'sd696;
		12'd2766: coeff = 10'sd695;
		12'd2767: coeff = 10'sd695;
		12'd2768: coeff = 10'sd694;
		12'd2769: coeff = 10'sd693;
		12'd2770: coeff = 10'sd692;
		12'd2771: coeff = 10'sd692;
		12'd2772: coeff = 10'sd691;
		12'd2773: coeff = 10'sd690;
		12'd2774: coeff = 10'sd689;
		12'd2775: coeff = 10'sd689;
		12'd2776: coeff = 10'sd688;
		12'd2777: coeff = 10'sd687;
		12'd2778: coeff = 10'sd686;
		12'd2779: coeff = 10'sd686;
		12'd2780: coeff = 10'sd685;
		12'd2781: coeff = 10'sd684;
		12'd2782: coeff = 10'sd683;
		12'd2783: coeff = 10'sd683;
		12'd2784: coeff = 10'sd682;
		12'd2785: coeff = 10'sd681;
		12'd2786: coeff = 10'sd680;
		12'd2787: coeff = 10'sd680;
		12'd2788: coeff = 10'sd679;
		12'd2789: coeff = 10'sd678;
		12'd2790: coeff = 10'sd677;
		12'd2791: coeff = 10'sd677;
		12'd2792: coeff = 10'sd676;
		12'd2793: coeff = 10'sd675;
		12'd2794: coeff = 10'sd674;
		12'd2795: coeff = 10'sd674;
		12'd2796: coeff = 10'sd673;
		12'd2797: coeff = 10'sd672;
		12'd2798: coeff = 10'sd671;
		12'd2799: coeff = 10'sd670;
		12'd2800: coeff = 10'sd670;
		12'd2801: coeff = 10'sd669;
		12'd2802: coeff = 10'sd668;
		12'd2803: coeff = 10'sd667;
		12'd2804: coeff = 10'sd667;
		12'd2805: coeff = 10'sd666;
		12'd2806: coeff = 10'sd665;
		12'd2807: coeff = 10'sd664;
		12'd2808: coeff = 10'sd664;
		12'd2809: coeff = 10'sd663;
		12'd2810: coeff = 10'sd662;
		12'd2811: coeff = 10'sd661;
		12'd2812: coeff = 10'sd660;
		12'd2813: coeff = 10'sd660;
		12'd2814: coeff = 10'sd659;
		12'd2815: coeff = 10'sd658;
		12'd2816: coeff = 10'sd657;
		12'd2817: coeff = 10'sd657;
		12'd2818: coeff = 10'sd656;
		12'd2819: coeff = 10'sd655;
		12'd2820: coeff = 10'sd654;
		12'd2821: coeff = 10'sd654;
		12'd2822: coeff = 10'sd653;
		12'd2823: coeff = 10'sd652;
		12'd2824: coeff = 10'sd651;
		12'd2825: coeff = 10'sd650;
		12'd2826: coeff = 10'sd650;
		12'd2827: coeff = 10'sd649;
		12'd2828: coeff = 10'sd648;
		12'd2829: coeff = 10'sd647;
		12'd2830: coeff = 10'sd647;
		12'd2831: coeff = 10'sd646;
		12'd2832: coeff = 10'sd645;
		12'd2833: coeff = 10'sd644;
		12'd2834: coeff = 10'sd643;
		12'd2835: coeff = 10'sd643;
		12'd2836: coeff = 10'sd642;
		12'd2837: coeff = 10'sd641;
		12'd2838: coeff = 10'sd640;
		12'd2839: coeff = 10'sd640;
		12'd2840: coeff = 10'sd639;
		12'd2841: coeff = 10'sd638;
		12'd2842: coeff = 10'sd637;
		12'd2843: coeff = 10'sd636;
		12'd2844: coeff = 10'sd636;
		12'd2845: coeff = 10'sd635;
		12'd2846: coeff = 10'sd634;
		12'd2847: coeff = 10'sd633;
		12'd2848: coeff = 10'sd633;
		12'd2849: coeff = 10'sd632;
		12'd2850: coeff = 10'sd631;
		12'd2851: coeff = 10'sd630;
		12'd2852: coeff = 10'sd629;
		12'd2853: coeff = 10'sd629;
		12'd2854: coeff = 10'sd628;
		12'd2855: coeff = 10'sd627;
		12'd2856: coeff = 10'sd626;
		12'd2857: coeff = 10'sd625;
		12'd2858: coeff = 10'sd625;
		12'd2859: coeff = 10'sd624;
		12'd2860: coeff = 10'sd623;
		12'd2861: coeff = 10'sd622;
		12'd2862: coeff = 10'sd622;
		12'd2863: coeff = 10'sd621;
		12'd2864: coeff = 10'sd620;
		12'd2865: coeff = 10'sd619;
		12'd2866: coeff = 10'sd618;
		12'd2867: coeff = 10'sd618;
		12'd2868: coeff = 10'sd617;
		12'd2869: coeff = 10'sd616;
		12'd2870: coeff = 10'sd615;
		12'd2871: coeff = 10'sd614;
		12'd2872: coeff = 10'sd614;
		12'd2873: coeff = 10'sd613;
		12'd2874: coeff = 10'sd612;
		12'd2875: coeff = 10'sd611;
		12'd2876: coeff = 10'sd611;
		12'd2877: coeff = 10'sd610;
		12'd2878: coeff = 10'sd609;
		12'd2879: coeff = 10'sd608;
		12'd2880: coeff = 10'sd607;
		12'd2881: coeff = 10'sd607;
		12'd2882: coeff = 10'sd606;
		12'd2883: coeff = 10'sd605;
		12'd2884: coeff = 10'sd604;
		12'd2885: coeff = 10'sd603;
		12'd2886: coeff = 10'sd603;
		12'd2887: coeff = 10'sd602;
		12'd2888: coeff = 10'sd601;
		12'd2889: coeff = 10'sd600;
		12'd2890: coeff = 10'sd599;
		12'd2891: coeff = 10'sd599;
		12'd2892: coeff = 10'sd598;
		12'd2893: coeff = 10'sd597;
		12'd2894: coeff = 10'sd596;
		12'd2895: coeff = 10'sd595;
		12'd2896: coeff = 10'sd595;
		12'd2897: coeff = 10'sd594;
		12'd2898: coeff = 10'sd593;
		12'd2899: coeff = 10'sd592;
		12'd2900: coeff = 10'sd592;
		12'd2901: coeff = 10'sd591;
		12'd2902: coeff = 10'sd590;
		12'd2903: coeff = 10'sd589;
		12'd2904: coeff = 10'sd588;
		12'd2905: coeff = 10'sd588;
		12'd2906: coeff = 10'sd587;
		12'd2907: coeff = 10'sd586;
		12'd2908: coeff = 10'sd585;
		12'd2909: coeff = 10'sd584;
		12'd2910: coeff = 10'sd584;
		12'd2911: coeff = 10'sd583;
		12'd2912: coeff = 10'sd582;
		12'd2913: coeff = 10'sd581;
		12'd2914: coeff = 10'sd580;
		12'd2915: coeff = 10'sd580;
		12'd2916: coeff = 10'sd579;
		12'd2917: coeff = 10'sd578;
		12'd2918: coeff = 10'sd577;
		12'd2919: coeff = 10'sd576;
		12'd2920: coeff = 10'sd576;
		12'd2921: coeff = 10'sd575;
		12'd2922: coeff = 10'sd574;
		12'd2923: coeff = 10'sd573;
		12'd2924: coeff = 10'sd572;
		12'd2925: coeff = 10'sd572;
		12'd2926: coeff = 10'sd571;
		12'd2927: coeff = 10'sd570;
		12'd2928: coeff = 10'sd569;
		12'd2929: coeff = 10'sd568;
		12'd2930: coeff = 10'sd568;
		12'd2931: coeff = 10'sd567;
		12'd2932: coeff = 10'sd566;
		12'd2933: coeff = 10'sd565;
		12'd2934: coeff = 10'sd564;
		12'd2935: coeff = 10'sd564;
		12'd2936: coeff = 10'sd563;
		12'd2937: coeff = 10'sd562;
		12'd2938: coeff = 10'sd561;
		12'd2939: coeff = 10'sd560;
		12'd2940: coeff = 10'sd560;
		12'd2941: coeff = 10'sd559;
		12'd2942: coeff = 10'sd558;
		12'd2943: coeff = 10'sd557;
		12'd2944: coeff = 10'sd556;
		12'd2945: coeff = 10'sd556;
		12'd2946: coeff = 10'sd555;
		12'd2947: coeff = 10'sd554;
		12'd2948: coeff = 10'sd553;
		12'd2949: coeff = 10'sd552;
		12'd2950: coeff = 10'sd552;
		12'd2951: coeff = 10'sd551;
		12'd2952: coeff = 10'sd550;
		12'd2953: coeff = 10'sd549;
		12'd2954: coeff = 10'sd548;
		12'd2955: coeff = 10'sd548;
		12'd2956: coeff = 10'sd547;
		12'd2957: coeff = 10'sd546;
		12'd2958: coeff = 10'sd545;
		12'd2959: coeff = 10'sd544;
		12'd2960: coeff = 10'sd544;
		12'd2961: coeff = 10'sd543;
		12'd2962: coeff = 10'sd542;
		12'd2963: coeff = 10'sd541;
		12'd2964: coeff = 10'sd540;
		12'd2965: coeff = 10'sd540;
		12'd2966: coeff = 10'sd539;
		12'd2967: coeff = 10'sd538;
		12'd2968: coeff = 10'sd537;
		12'd2969: coeff = 10'sd536;
		12'd2970: coeff = 10'sd536;
		12'd2971: coeff = 10'sd535;
		12'd2972: coeff = 10'sd534;
		12'd2973: coeff = 10'sd533;
		12'd2974: coeff = 10'sd532;
		12'd2975: coeff = 10'sd532;
		12'd2976: coeff = 10'sd531;
		12'd2977: coeff = 10'sd530;
		12'd2978: coeff = 10'sd529;
		12'd2979: coeff = 10'sd528;
		12'd2980: coeff = 10'sd527;
		12'd2981: coeff = 10'sd527;
		12'd2982: coeff = 10'sd526;
		12'd2983: coeff = 10'sd525;
		12'd2984: coeff = 10'sd524;
		12'd2985: coeff = 10'sd523;
		12'd2986: coeff = 10'sd523;
		12'd2987: coeff = 10'sd522;
		12'd2988: coeff = 10'sd521;
		12'd2989: coeff = 10'sd520;
		12'd2990: coeff = 10'sd519;
		12'd2991: coeff = 10'sd519;
		12'd2992: coeff = 10'sd518;
		12'd2993: coeff = 10'sd517;
		12'd2994: coeff = 10'sd516;
		12'd2995: coeff = 10'sd515;
		12'd2996: coeff = 10'sd515;
		12'd2997: coeff = 10'sd514;
		12'd2998: coeff = 10'sd513;
		12'd2999: coeff = 10'sd512;
		12'd3000: coeff = 10'sd511;
		12'd3001: coeff = 10'sd511;
		12'd3002: coeff = 10'sd510;
		12'd3003: coeff = 10'sd509;
		12'd3004: coeff = 10'sd508;
		12'd3005: coeff = 10'sd507;
		12'd3006: coeff = 10'sd507;
		12'd3007: coeff = 10'sd506;
		12'd3008: coeff = 10'sd505;
		12'd3009: coeff = 10'sd504;
		12'd3010: coeff = 10'sd503;
		12'd3011: coeff = 10'sd503;
		12'd3012: coeff = 10'sd502;
		12'd3013: coeff = 10'sd501;
		12'd3014: coeff = 10'sd500;
		12'd3015: coeff = 10'sd499;
		12'd3016: coeff = 10'sd499;
		12'd3017: coeff = 10'sd498;
		12'd3018: coeff = 10'sd497;
		12'd3019: coeff = 10'sd496;
		12'd3020: coeff = 10'sd495;
		12'd3021: coeff = 10'sd495;
		12'd3022: coeff = 10'sd494;
		12'd3023: coeff = 10'sd493;
		12'd3024: coeff = 10'sd492;
		12'd3025: coeff = 10'sd491;
		12'd3026: coeff = 10'sd490;
		12'd3027: coeff = 10'sd490;
		12'd3028: coeff = 10'sd489;
		12'd3029: coeff = 10'sd488;
		12'd3030: coeff = 10'sd487;
		12'd3031: coeff = 10'sd486;
		12'd3032: coeff = 10'sd486;
		12'd3033: coeff = 10'sd485;
		12'd3034: coeff = 10'sd484;
		12'd3035: coeff = 10'sd483;
		12'd3036: coeff = 10'sd482;
		12'd3037: coeff = 10'sd482;
		12'd3038: coeff = 10'sd481;
		12'd3039: coeff = 10'sd480;
		12'd3040: coeff = 10'sd479;
		12'd3041: coeff = 10'sd478;
		12'd3042: coeff = 10'sd478;
		12'd3043: coeff = 10'sd477;
		12'd3044: coeff = 10'sd476;
		12'd3045: coeff = 10'sd475;
		12'd3046: coeff = 10'sd474;
		12'd3047: coeff = 10'sd474;
		12'd3048: coeff = 10'sd473;
		12'd3049: coeff = 10'sd472;
		12'd3050: coeff = 10'sd471;
		12'd3051: coeff = 10'sd470;
		12'd3052: coeff = 10'sd470;
		12'd3053: coeff = 10'sd469;
		12'd3054: coeff = 10'sd468;
		12'd3055: coeff = 10'sd467;
		12'd3056: coeff = 10'sd466;
		12'd3057: coeff = 10'sd466;
		12'd3058: coeff = 10'sd465;
		12'd3059: coeff = 10'sd464;
		12'd3060: coeff = 10'sd463;
		12'd3061: coeff = 10'sd462;
		12'd3062: coeff = 10'sd462;
		12'd3063: coeff = 10'sd461;
		12'd3064: coeff = 10'sd460;
		12'd3065: coeff = 10'sd459;
		12'd3066: coeff = 10'sd458;
		12'd3067: coeff = 10'sd458;
		12'd3068: coeff = 10'sd457;
		12'd3069: coeff = 10'sd456;
		12'd3070: coeff = 10'sd455;
		12'd3071: coeff = 10'sd454;
		12'd3072: coeff = 10'sd454;
		12'd3073: coeff = 10'sd453;
		12'd3074: coeff = 10'sd452;
		12'd3075: coeff = 10'sd451;
		12'd3076: coeff = 10'sd450;
		12'd3077: coeff = 10'sd450;
		12'd3078: coeff = 10'sd449;
		12'd3079: coeff = 10'sd448;
		12'd3080: coeff = 10'sd447;
		12'd3081: coeff = 10'sd446;
		12'd3082: coeff = 10'sd446;
		12'd3083: coeff = 10'sd445;
		12'd3084: coeff = 10'sd444;
		12'd3085: coeff = 10'sd443;
		12'd3086: coeff = 10'sd442;
		12'd3087: coeff = 10'sd442;
		12'd3088: coeff = 10'sd441;
		12'd3089: coeff = 10'sd440;
		12'd3090: coeff = 10'sd439;
		12'd3091: coeff = 10'sd438;
		12'd3092: coeff = 10'sd438;
		12'd3093: coeff = 10'sd437;
		12'd3094: coeff = 10'sd436;
		12'd3095: coeff = 10'sd435;
		12'd3096: coeff = 10'sd434;
		12'd3097: coeff = 10'sd434;
		12'd3098: coeff = 10'sd433;
		12'd3099: coeff = 10'sd432;
		12'd3100: coeff = 10'sd431;
		12'd3101: coeff = 10'sd430;
		12'd3102: coeff = 10'sd430;
		12'd3103: coeff = 10'sd429;
		12'd3104: coeff = 10'sd428;
		12'd3105: coeff = 10'sd427;
		12'd3106: coeff = 10'sd427;
		12'd3107: coeff = 10'sd426;
		12'd3108: coeff = 10'sd425;
		12'd3109: coeff = 10'sd424;
		12'd3110: coeff = 10'sd423;
		12'd3111: coeff = 10'sd423;
		12'd3112: coeff = 10'sd422;
		12'd3113: coeff = 10'sd421;
		12'd3114: coeff = 10'sd420;
		12'd3115: coeff = 10'sd419;
		12'd3116: coeff = 10'sd419;
		12'd3117: coeff = 10'sd418;
		12'd3118: coeff = 10'sd417;
		12'd3119: coeff = 10'sd416;
		12'd3120: coeff = 10'sd415;
		12'd3121: coeff = 10'sd415;
		12'd3122: coeff = 10'sd414;
		12'd3123: coeff = 10'sd413;
		12'd3124: coeff = 10'sd412;
		12'd3125: coeff = 10'sd411;
		12'd3126: coeff = 10'sd411;
		12'd3127: coeff = 10'sd410;
		12'd3128: coeff = 10'sd409;
		12'd3129: coeff = 10'sd408;
		12'd3130: coeff = 10'sd408;
		12'd3131: coeff = 10'sd407;
		12'd3132: coeff = 10'sd406;
		12'd3133: coeff = 10'sd405;
		12'd3134: coeff = 10'sd404;
		12'd3135: coeff = 10'sd404;
		12'd3136: coeff = 10'sd403;
		12'd3137: coeff = 10'sd402;
		12'd3138: coeff = 10'sd401;
		12'd3139: coeff = 10'sd400;
		12'd3140: coeff = 10'sd400;
		12'd3141: coeff = 10'sd399;
		12'd3142: coeff = 10'sd398;
		12'd3143: coeff = 10'sd397;
		12'd3144: coeff = 10'sd397;
		12'd3145: coeff = 10'sd396;
		12'd3146: coeff = 10'sd395;
		12'd3147: coeff = 10'sd394;
		12'd3148: coeff = 10'sd393;
		12'd3149: coeff = 10'sd393;
		12'd3150: coeff = 10'sd392;
		12'd3151: coeff = 10'sd391;
		12'd3152: coeff = 10'sd390;
		12'd3153: coeff = 10'sd390;
		12'd3154: coeff = 10'sd389;
		12'd3155: coeff = 10'sd388;
		12'd3156: coeff = 10'sd387;
		12'd3157: coeff = 10'sd386;
		12'd3158: coeff = 10'sd386;
		12'd3159: coeff = 10'sd385;
		12'd3160: coeff = 10'sd384;
		12'd3161: coeff = 10'sd383;
		12'd3162: coeff = 10'sd382;
		12'd3163: coeff = 10'sd382;
		12'd3164: coeff = 10'sd381;
		12'd3165: coeff = 10'sd380;
		12'd3166: coeff = 10'sd379;
		12'd3167: coeff = 10'sd379;
		12'd3168: coeff = 10'sd378;
		12'd3169: coeff = 10'sd377;
		12'd3170: coeff = 10'sd376;
		12'd3171: coeff = 10'sd376;
		12'd3172: coeff = 10'sd375;
		12'd3173: coeff = 10'sd374;
		12'd3174: coeff = 10'sd373;
		12'd3175: coeff = 10'sd372;
		12'd3176: coeff = 10'sd372;
		12'd3177: coeff = 10'sd371;
		12'd3178: coeff = 10'sd370;
		12'd3179: coeff = 10'sd369;
		12'd3180: coeff = 10'sd369;
		12'd3181: coeff = 10'sd368;
		12'd3182: coeff = 10'sd367;
		12'd3183: coeff = 10'sd366;
		12'd3184: coeff = 10'sd365;
		12'd3185: coeff = 10'sd365;
		12'd3186: coeff = 10'sd364;
		12'd3187: coeff = 10'sd363;
		12'd3188: coeff = 10'sd362;
		12'd3189: coeff = 10'sd362;
		12'd3190: coeff = 10'sd361;
		12'd3191: coeff = 10'sd360;
		12'd3192: coeff = 10'sd359;
		12'd3193: coeff = 10'sd359;
		12'd3194: coeff = 10'sd358;
		12'd3195: coeff = 10'sd357;
		12'd3196: coeff = 10'sd356;
		12'd3197: coeff = 10'sd355;
		12'd3198: coeff = 10'sd355;
		12'd3199: coeff = 10'sd354;
		12'd3200: coeff = 10'sd353;
		12'd3201: coeff = 10'sd352;
		12'd3202: coeff = 10'sd352;
		12'd3203: coeff = 10'sd351;
		12'd3204: coeff = 10'sd350;
		12'd3205: coeff = 10'sd349;
		12'd3206: coeff = 10'sd349;
		12'd3207: coeff = 10'sd348;
		12'd3208: coeff = 10'sd347;
		12'd3209: coeff = 10'sd346;
		12'd3210: coeff = 10'sd346;
		12'd3211: coeff = 10'sd345;
		12'd3212: coeff = 10'sd344;
		12'd3213: coeff = 10'sd343;
		12'd3214: coeff = 10'sd343;
		12'd3215: coeff = 10'sd342;
		12'd3216: coeff = 10'sd341;
		12'd3217: coeff = 10'sd340;
		12'd3218: coeff = 10'sd339;
		12'd3219: coeff = 10'sd339;
		12'd3220: coeff = 10'sd338;
		12'd3221: coeff = 10'sd337;
		12'd3222: coeff = 10'sd336;
		12'd3223: coeff = 10'sd336;
		12'd3224: coeff = 10'sd335;
		12'd3225: coeff = 10'sd334;
		12'd3226: coeff = 10'sd333;
		12'd3227: coeff = 10'sd333;
		12'd3228: coeff = 10'sd332;
		12'd3229: coeff = 10'sd331;
		12'd3230: coeff = 10'sd330;
		12'd3231: coeff = 10'sd330;
		12'd3232: coeff = 10'sd329;
		12'd3233: coeff = 10'sd328;
		12'd3234: coeff = 10'sd327;
		12'd3235: coeff = 10'sd327;
		12'd3236: coeff = 10'sd326;
		12'd3237: coeff = 10'sd325;
		12'd3238: coeff = 10'sd324;
		12'd3239: coeff = 10'sd324;
		12'd3240: coeff = 10'sd323;
		12'd3241: coeff = 10'sd322;
		12'd3242: coeff = 10'sd321;
		12'd3243: coeff = 10'sd321;
		12'd3244: coeff = 10'sd320;
		12'd3245: coeff = 10'sd319;
		12'd3246: coeff = 10'sd318;
		12'd3247: coeff = 10'sd318;
		12'd3248: coeff = 10'sd317;
		12'd3249: coeff = 10'sd316;
		12'd3250: coeff = 10'sd315;
		12'd3251: coeff = 10'sd315;
		12'd3252: coeff = 10'sd314;
		12'd3253: coeff = 10'sd313;
		12'd3254: coeff = 10'sd312;
		12'd3255: coeff = 10'sd312;
		12'd3256: coeff = 10'sd311;
		12'd3257: coeff = 10'sd310;
		12'd3258: coeff = 10'sd310;
		12'd3259: coeff = 10'sd309;
		12'd3260: coeff = 10'sd308;
		12'd3261: coeff = 10'sd307;
		12'd3262: coeff = 10'sd307;
		12'd3263: coeff = 10'sd306;
		12'd3264: coeff = 10'sd305;
		12'd3265: coeff = 10'sd304;
		12'd3266: coeff = 10'sd304;
		12'd3267: coeff = 10'sd303;
		12'd3268: coeff = 10'sd302;
		12'd3269: coeff = 10'sd301;
		12'd3270: coeff = 10'sd301;
		12'd3271: coeff = 10'sd300;
		12'd3272: coeff = 10'sd299;
		12'd3273: coeff = 10'sd299;
		12'd3274: coeff = 10'sd298;
		12'd3275: coeff = 10'sd297;
		12'd3276: coeff = 10'sd296;
		12'd3277: coeff = 10'sd296;
		12'd3278: coeff = 10'sd295;
		12'd3279: coeff = 10'sd294;
		12'd3280: coeff = 10'sd293;
		12'd3281: coeff = 10'sd293;
		12'd3282: coeff = 10'sd292;
		12'd3283: coeff = 10'sd291;
		12'd3284: coeff = 10'sd290;
		12'd3285: coeff = 10'sd290;
		12'd3286: coeff = 10'sd289;
		12'd3287: coeff = 10'sd288;
		12'd3288: coeff = 10'sd288;
		12'd3289: coeff = 10'sd287;
		12'd3290: coeff = 10'sd286;
		12'd3291: coeff = 10'sd285;
		12'd3292: coeff = 10'sd285;
		12'd3293: coeff = 10'sd284;
		12'd3294: coeff = 10'sd283;
		12'd3295: coeff = 10'sd283;
		12'd3296: coeff = 10'sd282;
		12'd3297: coeff = 10'sd281;
		12'd3298: coeff = 10'sd280;
		12'd3299: coeff = 10'sd280;
		12'd3300: coeff = 10'sd279;
		12'd3301: coeff = 10'sd278;
		12'd3302: coeff = 10'sd278;
		12'd3303: coeff = 10'sd277;
		12'd3304: coeff = 10'sd276;
		12'd3305: coeff = 10'sd275;
		12'd3306: coeff = 10'sd275;
		12'd3307: coeff = 10'sd274;
		12'd3308: coeff = 10'sd273;
		12'd3309: coeff = 10'sd273;
		12'd3310: coeff = 10'sd272;
		12'd3311: coeff = 10'sd271;
		12'd3312: coeff = 10'sd270;
		12'd3313: coeff = 10'sd270;
		12'd3314: coeff = 10'sd269;
		12'd3315: coeff = 10'sd268;
		12'd3316: coeff = 10'sd268;
		12'd3317: coeff = 10'sd267;
		12'd3318: coeff = 10'sd266;
		12'd3319: coeff = 10'sd265;
		12'd3320: coeff = 10'sd265;
		12'd3321: coeff = 10'sd264;
		12'd3322: coeff = 10'sd263;
		12'd3323: coeff = 10'sd263;
		12'd3324: coeff = 10'sd262;
		12'd3325: coeff = 10'sd261;
		12'd3326: coeff = 10'sd261;
		12'd3327: coeff = 10'sd260;
		12'd3328: coeff = 10'sd259;
		12'd3329: coeff = 10'sd258;
		12'd3330: coeff = 10'sd258;
		12'd3331: coeff = 10'sd257;
		12'd3332: coeff = 10'sd256;
		12'd3333: coeff = 10'sd256;
		12'd3334: coeff = 10'sd255;
		12'd3335: coeff = 10'sd254;
		12'd3336: coeff = 10'sd254;
		12'd3337: coeff = 10'sd253;
		12'd3338: coeff = 10'sd252;
		12'd3339: coeff = 10'sd251;
		12'd3340: coeff = 10'sd251;
		12'd3341: coeff = 10'sd250;
		12'd3342: coeff = 10'sd249;
		12'd3343: coeff = 10'sd249;
		12'd3344: coeff = 10'sd248;
		12'd3345: coeff = 10'sd247;
		12'd3346: coeff = 10'sd247;
		12'd3347: coeff = 10'sd246;
		12'd3348: coeff = 10'sd245;
		12'd3349: coeff = 10'sd245;
		12'd3350: coeff = 10'sd244;
		12'd3351: coeff = 10'sd243;
		12'd3352: coeff = 10'sd243;
		12'd3353: coeff = 10'sd242;
		12'd3354: coeff = 10'sd241;
		12'd3355: coeff = 10'sd240;
		12'd3356: coeff = 10'sd240;
		12'd3357: coeff = 10'sd239;
		12'd3358: coeff = 10'sd238;
		12'd3359: coeff = 10'sd238;
		12'd3360: coeff = 10'sd237;
		12'd3361: coeff = 10'sd236;
		12'd3362: coeff = 10'sd236;
		12'd3363: coeff = 10'sd235;
		12'd3364: coeff = 10'sd234;
		12'd3365: coeff = 10'sd234;
		12'd3366: coeff = 10'sd233;
		12'd3367: coeff = 10'sd232;
		12'd3368: coeff = 10'sd232;
		12'd3369: coeff = 10'sd231;
		12'd3370: coeff = 10'sd230;
		12'd3371: coeff = 10'sd230;
		12'd3372: coeff = 10'sd229;
		12'd3373: coeff = 10'sd228;
		12'd3374: coeff = 10'sd228;
		12'd3375: coeff = 10'sd227;
		12'd3376: coeff = 10'sd226;
		12'd3377: coeff = 10'sd226;
		12'd3378: coeff = 10'sd225;
		12'd3379: coeff = 10'sd224;
		12'd3380: coeff = 10'sd224;
		12'd3381: coeff = 10'sd223;
		12'd3382: coeff = 10'sd222;
		12'd3383: coeff = 10'sd222;
		12'd3384: coeff = 10'sd221;
		12'd3385: coeff = 10'sd220;
		12'd3386: coeff = 10'sd220;
		12'd3387: coeff = 10'sd219;
		12'd3388: coeff = 10'sd218;
		12'd3389: coeff = 10'sd218;
		12'd3390: coeff = 10'sd217;
		12'd3391: coeff = 10'sd216;
		12'd3392: coeff = 10'sd216;
		12'd3393: coeff = 10'sd215;
		12'd3394: coeff = 10'sd214;
		12'd3395: coeff = 10'sd214;
		12'd3396: coeff = 10'sd213;
		12'd3397: coeff = 10'sd212;
		12'd3398: coeff = 10'sd212;
		12'd3399: coeff = 10'sd211;
		12'd3400: coeff = 10'sd211;
		12'd3401: coeff = 10'sd210;
		12'd3402: coeff = 10'sd209;
		12'd3403: coeff = 10'sd209;
		12'd3404: coeff = 10'sd208;
		12'd3405: coeff = 10'sd207;
		12'd3406: coeff = 10'sd207;
		12'd3407: coeff = 10'sd206;
		12'd3408: coeff = 10'sd205;
		12'd3409: coeff = 10'sd205;
		12'd3410: coeff = 10'sd204;
		12'd3411: coeff = 10'sd203;
		12'd3412: coeff = 10'sd203;
		12'd3413: coeff = 10'sd202;
		12'd3414: coeff = 10'sd201;
		12'd3415: coeff = 10'sd201;
		12'd3416: coeff = 10'sd200;
		12'd3417: coeff = 10'sd200;
		12'd3418: coeff = 10'sd199;
		12'd3419: coeff = 10'sd198;
		12'd3420: coeff = 10'sd198;
		12'd3421: coeff = 10'sd197;
		12'd3422: coeff = 10'sd196;
		12'd3423: coeff = 10'sd196;
		12'd3424: coeff = 10'sd195;
		12'd3425: coeff = 10'sd194;
		12'd3426: coeff = 10'sd194;
		12'd3427: coeff = 10'sd193;
		12'd3428: coeff = 10'sd193;
		12'd3429: coeff = 10'sd192;
		12'd3430: coeff = 10'sd191;
		12'd3431: coeff = 10'sd191;
		12'd3432: coeff = 10'sd190;
		12'd3433: coeff = 10'sd189;
		12'd3434: coeff = 10'sd189;
		12'd3435: coeff = 10'sd188;
		12'd3436: coeff = 10'sd188;
		12'd3437: coeff = 10'sd187;
		12'd3438: coeff = 10'sd186;
		12'd3439: coeff = 10'sd186;
		12'd3440: coeff = 10'sd185;
		12'd3441: coeff = 10'sd184;
		12'd3442: coeff = 10'sd184;
		12'd3443: coeff = 10'sd183;
		12'd3444: coeff = 10'sd183;
		12'd3445: coeff = 10'sd182;
		12'd3446: coeff = 10'sd181;
		12'd3447: coeff = 10'sd181;
		12'd3448: coeff = 10'sd180;
		12'd3449: coeff = 10'sd180;
		12'd3450: coeff = 10'sd179;
		12'd3451: coeff = 10'sd178;
		12'd3452: coeff = 10'sd178;
		12'd3453: coeff = 10'sd177;
		12'd3454: coeff = 10'sd177;
		12'd3455: coeff = 10'sd176;
		12'd3456: coeff = 10'sd175;
		12'd3457: coeff = 10'sd175;
		12'd3458: coeff = 10'sd174;
		12'd3459: coeff = 10'sd173;
		12'd3460: coeff = 10'sd173;
		12'd3461: coeff = 10'sd172;
		12'd3462: coeff = 10'sd172;
		12'd3463: coeff = 10'sd171;
		12'd3464: coeff = 10'sd170;
		12'd3465: coeff = 10'sd170;
		12'd3466: coeff = 10'sd169;
		12'd3467: coeff = 10'sd169;
		12'd3468: coeff = 10'sd168;
		12'd3469: coeff = 10'sd167;
		12'd3470: coeff = 10'sd167;
		12'd3471: coeff = 10'sd166;
		12'd3472: coeff = 10'sd166;
		12'd3473: coeff = 10'sd165;
		12'd3474: coeff = 10'sd165;
		12'd3475: coeff = 10'sd164;
		12'd3476: coeff = 10'sd163;
		12'd3477: coeff = 10'sd163;
		12'd3478: coeff = 10'sd162;
		12'd3479: coeff = 10'sd162;
		12'd3480: coeff = 10'sd161;
		12'd3481: coeff = 10'sd160;
		12'd3482: coeff = 10'sd160;
		12'd3483: coeff = 10'sd159;
		12'd3484: coeff = 10'sd159;
		12'd3485: coeff = 10'sd158;
		12'd3486: coeff = 10'sd158;
		12'd3487: coeff = 10'sd157;
		12'd3488: coeff = 10'sd156;
		12'd3489: coeff = 10'sd156;
		12'd3490: coeff = 10'sd155;
		12'd3491: coeff = 10'sd155;
		12'd3492: coeff = 10'sd154;
		12'd3493: coeff = 10'sd153;
		12'd3494: coeff = 10'sd153;
		12'd3495: coeff = 10'sd152;
		12'd3496: coeff = 10'sd152;
		12'd3497: coeff = 10'sd151;
		12'd3498: coeff = 10'sd151;
		12'd3499: coeff = 10'sd150;
		12'd3500: coeff = 10'sd149;
		12'd3501: coeff = 10'sd149;
		12'd3502: coeff = 10'sd148;
		12'd3503: coeff = 10'sd148;
		12'd3504: coeff = 10'sd147;
		12'd3505: coeff = 10'sd147;
		12'd3506: coeff = 10'sd146;
		12'd3507: coeff = 10'sd146;
		12'd3508: coeff = 10'sd145;
		12'd3509: coeff = 10'sd144;
		12'd3510: coeff = 10'sd144;
		12'd3511: coeff = 10'sd143;
		12'd3512: coeff = 10'sd143;
		12'd3513: coeff = 10'sd142;
		12'd3514: coeff = 10'sd142;
		12'd3515: coeff = 10'sd141;
		12'd3516: coeff = 10'sd140;
		12'd3517: coeff = 10'sd140;
		12'd3518: coeff = 10'sd139;
		12'd3519: coeff = 10'sd139;
		12'd3520: coeff = 10'sd138;
		12'd3521: coeff = 10'sd138;
		12'd3522: coeff = 10'sd137;
		12'd3523: coeff = 10'sd137;
		12'd3524: coeff = 10'sd136;
		12'd3525: coeff = 10'sd136;
		12'd3526: coeff = 10'sd135;
		12'd3527: coeff = 10'sd134;
		12'd3528: coeff = 10'sd134;
		12'd3529: coeff = 10'sd133;
		12'd3530: coeff = 10'sd133;
		12'd3531: coeff = 10'sd132;
		12'd3532: coeff = 10'sd132;
		12'd3533: coeff = 10'sd131;
		12'd3534: coeff = 10'sd131;
		12'd3535: coeff = 10'sd130;
		12'd3536: coeff = 10'sd130;
		12'd3537: coeff = 10'sd129;
		12'd3538: coeff = 10'sd129;
		12'd3539: coeff = 10'sd128;
		12'd3540: coeff = 10'sd127;
		12'd3541: coeff = 10'sd127;
		12'd3542: coeff = 10'sd126;
		12'd3543: coeff = 10'sd126;
		12'd3544: coeff = 10'sd125;
		12'd3545: coeff = 10'sd125;
		12'd3546: coeff = 10'sd124;
		12'd3547: coeff = 10'sd124;
		12'd3548: coeff = 10'sd123;
		12'd3549: coeff = 10'sd123;
		12'd3550: coeff = 10'sd122;
		12'd3551: coeff = 10'sd122;
		12'd3552: coeff = 10'sd121;
		12'd3553: coeff = 10'sd121;
		12'd3554: coeff = 10'sd120;
		12'd3555: coeff = 10'sd120;
		12'd3556: coeff = 10'sd119;
		12'd3557: coeff = 10'sd119;
		12'd3558: coeff = 10'sd118;
		12'd3559: coeff = 10'sd118;
		12'd3560: coeff = 10'sd117;
		12'd3561: coeff = 10'sd117;
		12'd3562: coeff = 10'sd116;
		12'd3563: coeff = 10'sd116;
		12'd3564: coeff = 10'sd115;
		12'd3565: coeff = 10'sd114;
		12'd3566: coeff = 10'sd114;
		12'd3567: coeff = 10'sd113;
		12'd3568: coeff = 10'sd113;
		12'd3569: coeff = 10'sd112;
		12'd3570: coeff = 10'sd112;
		12'd3571: coeff = 10'sd111;
		12'd3572: coeff = 10'sd111;
		12'd3573: coeff = 10'sd110;
		12'd3574: coeff = 10'sd110;
		12'd3575: coeff = 10'sd109;
		12'd3576: coeff = 10'sd109;
		12'd3577: coeff = 10'sd108;
		12'd3578: coeff = 10'sd108;
		12'd3579: coeff = 10'sd107;
		12'd3580: coeff = 10'sd107;
		12'd3581: coeff = 10'sd107;
		12'd3582: coeff = 10'sd106;
		12'd3583: coeff = 10'sd106;
		12'd3584: coeff = 10'sd105;
		12'd3585: coeff = 10'sd105;
		12'd3586: coeff = 10'sd104;
		12'd3587: coeff = 10'sd104;
		12'd3588: coeff = 10'sd103;
		12'd3589: coeff = 10'sd103;
		12'd3590: coeff = 10'sd102;
		12'd3591: coeff = 10'sd102;
		12'd3592: coeff = 10'sd101;
		12'd3593: coeff = 10'sd101;
		12'd3594: coeff = 10'sd100;
		12'd3595: coeff = 10'sd100;
		12'd3596: coeff = 10'sd99;
		12'd3597: coeff = 10'sd99;
		12'd3598: coeff = 10'sd98;
		12'd3599: coeff = 10'sd98;
		12'd3600: coeff = 10'sd97;
		12'd3601: coeff = 10'sd97;
		12'd3602: coeff = 10'sd96;
		12'd3603: coeff = 10'sd96;
		12'd3604: coeff = 10'sd95;
		12'd3605: coeff = 10'sd95;
		12'd3606: coeff = 10'sd95;
		12'd3607: coeff = 10'sd94;
		12'd3608: coeff = 10'sd94;
		12'd3609: coeff = 10'sd93;
		12'd3610: coeff = 10'sd93;
		12'd3611: coeff = 10'sd92;
		12'd3612: coeff = 10'sd92;
		12'd3613: coeff = 10'sd91;
		12'd3614: coeff = 10'sd91;
		12'd3615: coeff = 10'sd90;
		12'd3616: coeff = 10'sd90;
		12'd3617: coeff = 10'sd89;
		12'd3618: coeff = 10'sd89;
		12'd3619: coeff = 10'sd89;
		12'd3620: coeff = 10'sd88;
		12'd3621: coeff = 10'sd88;
		12'd3622: coeff = 10'sd87;
		12'd3623: coeff = 10'sd87;
		12'd3624: coeff = 10'sd86;
		12'd3625: coeff = 10'sd86;
		12'd3626: coeff = 10'sd85;
		12'd3627: coeff = 10'sd85;
		12'd3628: coeff = 10'sd85;
		12'd3629: coeff = 10'sd84;
		12'd3630: coeff = 10'sd84;
		12'd3631: coeff = 10'sd83;
		12'd3632: coeff = 10'sd83;
		12'd3633: coeff = 10'sd82;
		12'd3634: coeff = 10'sd82;
		12'd3635: coeff = 10'sd81;
		12'd3636: coeff = 10'sd81;
		12'd3637: coeff = 10'sd81;
		12'd3638: coeff = 10'sd80;
		12'd3639: coeff = 10'sd80;
		12'd3640: coeff = 10'sd79;
		12'd3641: coeff = 10'sd79;
		12'd3642: coeff = 10'sd78;
		12'd3643: coeff = 10'sd78;
		12'd3644: coeff = 10'sd78;
		12'd3645: coeff = 10'sd77;
		12'd3646: coeff = 10'sd77;
		12'd3647: coeff = 10'sd76;
		12'd3648: coeff = 10'sd76;
		12'd3649: coeff = 10'sd75;
		12'd3650: coeff = 10'sd75;
		12'd3651: coeff = 10'sd75;
		12'd3652: coeff = 10'sd74;
		12'd3653: coeff = 10'sd74;
		12'd3654: coeff = 10'sd73;
		12'd3655: coeff = 10'sd73;
		12'd3656: coeff = 10'sd73;
		12'd3657: coeff = 10'sd72;
		12'd3658: coeff = 10'sd72;
		12'd3659: coeff = 10'sd71;
		12'd3660: coeff = 10'sd71;
		12'd3661: coeff = 10'sd71;
		12'd3662: coeff = 10'sd70;
		12'd3663: coeff = 10'sd70;
		12'd3664: coeff = 10'sd69;
		12'd3665: coeff = 10'sd69;
		12'd3666: coeff = 10'sd68;
		12'd3667: coeff = 10'sd68;
		12'd3668: coeff = 10'sd68;
		12'd3669: coeff = 10'sd67;
		12'd3670: coeff = 10'sd67;
		12'd3671: coeff = 10'sd66;
		12'd3672: coeff = 10'sd66;
		12'd3673: coeff = 10'sd66;
		12'd3674: coeff = 10'sd65;
		12'd3675: coeff = 10'sd65;
		12'd3676: coeff = 10'sd65;
		12'd3677: coeff = 10'sd64;
		12'd3678: coeff = 10'sd64;
		12'd3679: coeff = 10'sd63;
		12'd3680: coeff = 10'sd63;
		12'd3681: coeff = 10'sd63;
		12'd3682: coeff = 10'sd62;
		12'd3683: coeff = 10'sd62;
		12'd3684: coeff = 10'sd61;
		12'd3685: coeff = 10'sd61;
		12'd3686: coeff = 10'sd61;
		12'd3687: coeff = 10'sd60;
		12'd3688: coeff = 10'sd60;
		12'd3689: coeff = 10'sd60;
		12'd3690: coeff = 10'sd59;
		12'd3691: coeff = 10'sd59;
		12'd3692: coeff = 10'sd58;
		12'd3693: coeff = 10'sd58;
		12'd3694: coeff = 10'sd58;
		12'd3695: coeff = 10'sd57;
		12'd3696: coeff = 10'sd57;
		12'd3697: coeff = 10'sd57;
		12'd3698: coeff = 10'sd56;
		12'd3699: coeff = 10'sd56;
		12'd3700: coeff = 10'sd55;
		12'd3701: coeff = 10'sd55;
		12'd3702: coeff = 10'sd55;
		12'd3703: coeff = 10'sd54;
		12'd3704: coeff = 10'sd54;
		12'd3705: coeff = 10'sd54;
		12'd3706: coeff = 10'sd53;
		12'd3707: coeff = 10'sd53;
		12'd3708: coeff = 10'sd53;
		12'd3709: coeff = 10'sd52;
		12'd3710: coeff = 10'sd52;
		12'd3711: coeff = 10'sd52;
		12'd3712: coeff = 10'sd51;
		12'd3713: coeff = 10'sd51;
		12'd3714: coeff = 10'sd50;
		12'd3715: coeff = 10'sd50;
		12'd3716: coeff = 10'sd50;
		12'd3717: coeff = 10'sd49;
		12'd3718: coeff = 10'sd49;
		12'd3719: coeff = 10'sd49;
		12'd3720: coeff = 10'sd48;
		12'd3721: coeff = 10'sd48;
		12'd3722: coeff = 10'sd48;
		12'd3723: coeff = 10'sd47;
		12'd3724: coeff = 10'sd47;
		12'd3725: coeff = 10'sd47;
		12'd3726: coeff = 10'sd46;
		12'd3727: coeff = 10'sd46;
		12'd3728: coeff = 10'sd46;
		12'd3729: coeff = 10'sd45;
		12'd3730: coeff = 10'sd45;
		12'd3731: coeff = 10'sd45;
		12'd3732: coeff = 10'sd44;
		12'd3733: coeff = 10'sd44;
		12'd3734: coeff = 10'sd44;
		12'd3735: coeff = 10'sd43;
		12'd3736: coeff = 10'sd43;
		12'd3737: coeff = 10'sd43;
		12'd3738: coeff = 10'sd42;
		12'd3739: coeff = 10'sd42;
		12'd3740: coeff = 10'sd42;
		12'd3741: coeff = 10'sd41;
		12'd3742: coeff = 10'sd41;
		12'd3743: coeff = 10'sd41;
		12'd3744: coeff = 10'sd41;
		12'd3745: coeff = 10'sd40;
		12'd3746: coeff = 10'sd40;
		12'd3747: coeff = 10'sd40;
		12'd3748: coeff = 10'sd39;
		12'd3749: coeff = 10'sd39;
		12'd3750: coeff = 10'sd39;
		12'd3751: coeff = 10'sd38;
		12'd3752: coeff = 10'sd38;
		12'd3753: coeff = 10'sd38;
		12'd3754: coeff = 10'sd37;
		12'd3755: coeff = 10'sd37;
		12'd3756: coeff = 10'sd37;
		12'd3757: coeff = 10'sd37;
		12'd3758: coeff = 10'sd36;
		12'd3759: coeff = 10'sd36;
		12'd3760: coeff = 10'sd36;
		12'd3761: coeff = 10'sd35;
		12'd3762: coeff = 10'sd35;
		12'd3763: coeff = 10'sd35;
		12'd3764: coeff = 10'sd35;
		12'd3765: coeff = 10'sd34;
		12'd3766: coeff = 10'sd34;
		12'd3767: coeff = 10'sd34;
		12'd3768: coeff = 10'sd33;
		12'd3769: coeff = 10'sd33;
		12'd3770: coeff = 10'sd33;
		12'd3771: coeff = 10'sd33;
		12'd3772: coeff = 10'sd32;
		12'd3773: coeff = 10'sd32;
		12'd3774: coeff = 10'sd32;
		12'd3775: coeff = 10'sd31;
		12'd3776: coeff = 10'sd31;
		12'd3777: coeff = 10'sd31;
		12'd3778: coeff = 10'sd31;
		12'd3779: coeff = 10'sd30;
		12'd3780: coeff = 10'sd30;
		12'd3781: coeff = 10'sd30;
		12'd3782: coeff = 10'sd29;
		12'd3783: coeff = 10'sd29;
		12'd3784: coeff = 10'sd29;
		12'd3785: coeff = 10'sd29;
		12'd3786: coeff = 10'sd28;
		12'd3787: coeff = 10'sd28;
		12'd3788: coeff = 10'sd28;
		12'd3789: coeff = 10'sd28;
		12'd3790: coeff = 10'sd27;
		12'd3791: coeff = 10'sd27;
		12'd3792: coeff = 10'sd27;
		12'd3793: coeff = 10'sd27;
		12'd3794: coeff = 10'sd26;
		12'd3795: coeff = 10'sd26;
		12'd3796: coeff = 10'sd26;
		12'd3797: coeff = 10'sd26;
		12'd3798: coeff = 10'sd25;
		12'd3799: coeff = 10'sd25;
		12'd3800: coeff = 10'sd25;
		12'd3801: coeff = 10'sd25;
		12'd3802: coeff = 10'sd24;
		12'd3803: coeff = 10'sd24;
		12'd3804: coeff = 10'sd24;
		12'd3805: coeff = 10'sd24;
		12'd3806: coeff = 10'sd23;
		12'd3807: coeff = 10'sd23;
		12'd3808: coeff = 10'sd23;
		12'd3809: coeff = 10'sd23;
		12'd3810: coeff = 10'sd22;
		12'd3811: coeff = 10'sd22;
		12'd3812: coeff = 10'sd22;
		12'd3813: coeff = 10'sd22;
		12'd3814: coeff = 10'sd21;
		12'd3815: coeff = 10'sd21;
		12'd3816: coeff = 10'sd21;
		12'd3817: coeff = 10'sd21;
		12'd3818: coeff = 10'sd21;
		12'd3819: coeff = 10'sd20;
		12'd3820: coeff = 10'sd20;
		12'd3821: coeff = 10'sd20;
		12'd3822: coeff = 10'sd20;
		12'd3823: coeff = 10'sd19;
		12'd3824: coeff = 10'sd19;
		12'd3825: coeff = 10'sd19;
		12'd3826: coeff = 10'sd19;
		12'd3827: coeff = 10'sd19;
		12'd3828: coeff = 10'sd18;
		12'd3829: coeff = 10'sd18;
		12'd3830: coeff = 10'sd18;
		12'd3831: coeff = 10'sd18;
		12'd3832: coeff = 10'sd18;
		12'd3833: coeff = 10'sd17;
		12'd3834: coeff = 10'sd17;
		12'd3835: coeff = 10'sd17;
		12'd3836: coeff = 10'sd17;
		12'd3837: coeff = 10'sd16;
		12'd3838: coeff = 10'sd16;
		12'd3839: coeff = 10'sd16;
		12'd3840: coeff = 10'sd16;
		12'd3841: coeff = 10'sd16;
		12'd3842: coeff = 10'sd15;
		12'd3843: coeff = 10'sd15;
		12'd3844: coeff = 10'sd15;
		12'd3845: coeff = 10'sd15;
		12'd3846: coeff = 10'sd15;
		12'd3847: coeff = 10'sd15;
		12'd3848: coeff = 10'sd14;
		12'd3849: coeff = 10'sd14;
		12'd3850: coeff = 10'sd14;
		12'd3851: coeff = 10'sd14;
		12'd3852: coeff = 10'sd14;
		12'd3853: coeff = 10'sd13;
		12'd3854: coeff = 10'sd13;
		12'd3855: coeff = 10'sd13;
		12'd3856: coeff = 10'sd13;
		12'd3857: coeff = 10'sd13;
		12'd3858: coeff = 10'sd13;
		12'd3859: coeff = 10'sd12;
		12'd3860: coeff = 10'sd12;
		12'd3861: coeff = 10'sd12;
		12'd3862: coeff = 10'sd12;
		12'd3863: coeff = 10'sd12;
		12'd3864: coeff = 10'sd11;
		12'd3865: coeff = 10'sd11;
		12'd3866: coeff = 10'sd11;
		12'd3867: coeff = 10'sd11;
		12'd3868: coeff = 10'sd11;
		12'd3869: coeff = 10'sd11;
		12'd3870: coeff = 10'sd10;
		12'd3871: coeff = 10'sd10;
		12'd3872: coeff = 10'sd10;
		12'd3873: coeff = 10'sd10;
		12'd3874: coeff = 10'sd10;
		12'd3875: coeff = 10'sd10;
		12'd3876: coeff = 10'sd10;
		12'd3877: coeff = 10'sd9;
		12'd3878: coeff = 10'sd9;
		12'd3879: coeff = 10'sd9;
		12'd3880: coeff = 10'sd9;
		12'd3881: coeff = 10'sd9;
		12'd3882: coeff = 10'sd9;
		12'd3883: coeff = 10'sd8;
		12'd3884: coeff = 10'sd8;
		12'd3885: coeff = 10'sd8;
		12'd3886: coeff = 10'sd8;
		12'd3887: coeff = 10'sd8;
		12'd3888: coeff = 10'sd8;
		12'd3889: coeff = 10'sd8;
		12'd3890: coeff = 10'sd7;
		12'd3891: coeff = 10'sd7;
		12'd3892: coeff = 10'sd7;
		12'd3893: coeff = 10'sd7;
		12'd3894: coeff = 10'sd7;
		12'd3895: coeff = 10'sd7;
		12'd3896: coeff = 10'sd7;
		12'd3897: coeff = 10'sd7;
		12'd3898: coeff = 10'sd6;
		12'd3899: coeff = 10'sd6;
		12'd3900: coeff = 10'sd6;
		12'd3901: coeff = 10'sd6;
		12'd3902: coeff = 10'sd6;
		12'd3903: coeff = 10'sd6;
		12'd3904: coeff = 10'sd6;
		12'd3905: coeff = 10'sd6;
		12'd3906: coeff = 10'sd5;
		12'd3907: coeff = 10'sd5;
		12'd3908: coeff = 10'sd5;
		12'd3909: coeff = 10'sd5;
		12'd3910: coeff = 10'sd5;
		12'd3911: coeff = 10'sd5;
		12'd3912: coeff = 10'sd5;
		12'd3913: coeff = 10'sd5;
		12'd3914: coeff = 10'sd5;
		12'd3915: coeff = 10'sd4;
		12'd3916: coeff = 10'sd4;
		12'd3917: coeff = 10'sd4;
		12'd3918: coeff = 10'sd4;
		12'd3919: coeff = 10'sd4;
		12'd3920: coeff = 10'sd4;
		12'd3921: coeff = 10'sd4;
		12'd3922: coeff = 10'sd4;
		12'd3923: coeff = 10'sd4;
		12'd3924: coeff = 10'sd4;
		12'd3925: coeff = 10'sd3;
		12'd3926: coeff = 10'sd3;
		12'd3927: coeff = 10'sd3;
		12'd3928: coeff = 10'sd3;
		12'd3929: coeff = 10'sd3;
		12'd3930: coeff = 10'sd3;
		12'd3931: coeff = 10'sd3;
		12'd3932: coeff = 10'sd3;
		12'd3933: coeff = 10'sd3;
		12'd3934: coeff = 10'sd3;
		12'd3935: coeff = 10'sd3;
		12'd3936: coeff = 10'sd3;
		12'd3937: coeff = 10'sd2;
		12'd3938: coeff = 10'sd2;
		12'd3939: coeff = 10'sd2;
		12'd3940: coeff = 10'sd2;
		12'd3941: coeff = 10'sd2;
		12'd3942: coeff = 10'sd2;
		12'd3943: coeff = 10'sd2;
		12'd3944: coeff = 10'sd2;
		12'd3945: coeff = 10'sd2;
		12'd3946: coeff = 10'sd2;
		12'd3947: coeff = 10'sd2;
		12'd3948: coeff = 10'sd2;
		12'd3949: coeff = 10'sd2;
		12'd3950: coeff = 10'sd2;
		12'd3951: coeff = 10'sd1;
		12'd3952: coeff = 10'sd1;
		12'd3953: coeff = 10'sd1;
		12'd3954: coeff = 10'sd1;
		12'd3955: coeff = 10'sd1;
		12'd3956: coeff = 10'sd1;
		12'd3957: coeff = 10'sd1;
		12'd3958: coeff = 10'sd1;
		12'd3959: coeff = 10'sd1;
		12'd3960: coeff = 10'sd1;
		12'd3961: coeff = 10'sd1;
		12'd3962: coeff = 10'sd1;
		12'd3963: coeff = 10'sd1;
		12'd3964: coeff = 10'sd1;
		12'd3965: coeff = 10'sd1;
		12'd3966: coeff = 10'sd1;
		12'd3967: coeff = 10'sd1;
		12'd3968: coeff = 10'sd1;
		12'd3969: coeff = 10'sd1;
		12'd3970: coeff = 10'sd1;
		12'd3971: coeff = 10'sd0;
		12'd3972: coeff = 10'sd0;
		12'd3973: coeff = 10'sd0;
		12'd3974: coeff = 10'sd0;
		12'd3975: coeff = 10'sd0;
		12'd3976: coeff = 10'sd0;
		12'd3977: coeff = 10'sd0;
		12'd3978: coeff = 10'sd0;
		12'd3979: coeff = 10'sd0;
		12'd3980: coeff = 10'sd0;
		12'd3981: coeff = 10'sd0;
		12'd3982: coeff = 10'sd0;
		12'd3983: coeff = 10'sd0;
		12'd3984: coeff = 10'sd0;
		12'd3985: coeff = 10'sd0;
		12'd3986: coeff = 10'sd0;
		12'd3987: coeff = 10'sd0;
		12'd3988: coeff = 10'sd0;
		12'd3989: coeff = 10'sd0;
		12'd3990: coeff = 10'sd0;
		12'd3991: coeff = 10'sd0;
		12'd3992: coeff = 10'sd0;
		12'd3993: coeff = 10'sd0;
		12'd3994: coeff = 10'sd0;
		12'd3995: coeff = 10'sd0;
		12'd3996: coeff = 10'sd0;
		12'd3997: coeff = 10'sd0;
		12'd3998: coeff = 10'sd0;
		12'd3999: coeff = 10'sd0;
		endcase
endmodule
